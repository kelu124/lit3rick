interface mi_if;
    bit clk;
    bit reset;

    bit top_turn2;
    bit BUT_USER;
    bit BUT_TRIG;
endinterface