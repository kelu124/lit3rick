module chip (io_12_31_1, io_13_0_1, io_13_31_0, io_13_31_1, io_15_0_0, io_16_0_0, io_16_31_0, io_16_31_1, io_17_0_0, io_17_31_0, io_18_0_0, io_18_0_1, io_18_31_0, io_18_31_1, io_19_0_0, io_19_0_1, io_21_0_1, io_22_0_1, io_23_0_0, io_23_0_1, io_4_31_0, io_5_0_0, io_5_31_0, io_6_0_0, io_6_0_1, io_6_31_0, io_7_0_0, io_8_0_0, io_8_31_0, io_8_31_1, io_9_0_0, io_9_0_1);
  wire net_5;
  wire net_6;
  wire net_8;
  wire net_9;
  wire net_10;
  wire net_12;
  wire net_103;
  wire net_106;
  wire net_107;
  wire net_108;
  wire net_117;
  wire net_118;
  wire net_119;
  wire net_120;
  wire net_121;
  wire net_122;
  wire net_123;
  wire net_250;
  wire net_292;
  wire net_451;
  wire net_452;
  wire net_453;
  wire net_454;
  wire net_455;
  wire net_456;
  wire net_457;
  wire net_458;
  wire net_523;
  wire net_571;
  wire net_679;
  wire net_680;
  wire net_681;
  wire net_682;
  wire net_683;
  wire net_684;
  wire net_685;
  wire net_761;
  wire net_788;
  wire net_798;
  wire net_804;
  wire net_811;
  wire net_905;
  wire net_906;
  wire net_907;
  wire net_908;
  wire net_909;
  wire net_910;
  wire net_911;
  wire net_912;
  wire net_1017;
  wire net_1019;
  wire net_1023;
  wire net_1027;
  wire net_1031;
  wire net_1037;
  wire net_1098;
  wire net_1099;
  wire net_1100;
  wire net_1101;
  wire net_1102;
  wire net_1103;
  wire net_1104;
  wire net_1105;
  wire net_1131;
  wire net_1133;
  wire net_1134;
  wire net_1135;
  wire net_1136;
  wire net_1178;
  wire net_1181;
  wire net_1184;
  wire net_1195;
  wire net_1199;
  wire net_1201;
  wire net_1206;
  wire net_1210;
  wire net_1223;
  wire net_1224;
  wire net_1225;
  wire net_1227;
  wire net_1228;
  wire net_1232;
  wire net_1233;
  wire net_1235;
  wire net_1236;
  wire net_1257;
  wire net_1258;
  wire net_1259;
  wire net_1262;
  wire net_1264;
  wire net_1267;
  wire net_1268;
  wire net_1272;
  wire net_1274;
  wire net_1275;
  wire net_1276;
  wire net_1278;
  wire net_1279;
  wire net_1280;
  wire net_1281;
  wire net_1285;
  wire net_1287;
  wire net_1288;
  wire net_1289;
  wire net_1290;
  wire net_1291;
  wire net_1292;
  wire net_1293;
  wire net_1294;
  wire net_1295;
  wire net_1296;
  wire net_1297;
  wire net_1298;
  wire net_1299;
  wire net_1300;
  wire net_1301;
  wire net_1302;
  wire net_1304;
  wire net_1305;
  wire net_1306;
  wire net_1307;
  wire net_1308;
  wire net_1309;
  wire net_1310;
  wire net_1311;
  wire net_1337;
  wire net_1384;
  wire net_1386;
  wire net_1418;
  wire net_1423;
  wire net_1430;
  wire net_1436;
  wire net_1440;
  wire net_1447;
  wire net_1461;
  wire net_1464;
  wire net_1471;
  wire net_1474;
  wire net_1476;
  wire net_1478;
  wire net_1479;
  wire net_1483;
  wire net_1484;
  wire net_1485;
  wire net_1486;
  wire net_1487;
  wire net_1488;
  wire net_1489;
  wire net_1490;
  wire net_1491;
  wire net_1493;
  wire net_1494;
  wire net_1495;
  wire net_1496;
  wire net_1497;
  wire net_1498;
  wire net_1499;
  wire net_1500;
  wire net_1501;
  wire net_1502;
  wire net_1503;
  wire net_1504;
  wire net_1505;
  wire net_1506;
  wire net_1507;
  wire net_1508;
  wire net_1512;
  wire net_1513;
  wire net_1514;
  wire net_1515;
  wire net_1516;
  wire net_1517;
  wire net_1518;
  wire net_1519;
  wire net_1544;
  wire net_1545;
  wire net_1546;
  wire net_1547;
  wire net_1548;
  wire net_1549;
  wire net_1550;
  wire net_1551;
  wire net_1555;
  wire net_1594;
  wire net_1598;
  wire net_1618;
  wire net_1636;
  wire net_1645;
  wire net_1647;
  wire net_1656;
  wire net_1658;
  wire net_1721;
  wire net_1722;
  wire net_1723;
  wire net_1724;
  wire net_1725;
  wire net_1726;
  wire net_1727;
  wire net_1753;
  wire net_1754;
  wire net_1755;
  wire net_1756;
  wire net_1757;
  wire net_1758;
  wire net_1759;
  wire net_1760;
  wire net_1764;
  wire net_1801;
  wire net_1805;
  wire net_1814;
  wire net_1850;
  wire net_1851;
  wire net_1853;
  wire net_1856;
  wire net_1858;
  wire net_1860;
  wire net_1965;
  wire net_1966;
  wire net_1967;
  wire net_1968;
  wire net_1969;
  wire net_1970;
  wire net_1971;
  wire net_1972;
  wire net_1991;
  wire net_1992;
  wire net_2002;
  wire net_2012;
  wire net_2071;
  wire net_2076;
  wire net_2078;
  wire net_2086;
  wire net_2088;
  wire net_2158;
  wire net_2159;
  wire net_2160;
  wire net_2161;
  wire net_2162;
  wire net_2163;
  wire net_2164;
  wire net_2165;
  wire net_2190;
  wire net_2191;
  wire net_2192;
  wire net_2193;
  wire net_2194;
  wire net_2195;
  wire net_2196;
  wire net_2197;
  wire net_2200;
  wire net_2239;
  wire net_2248;
  wire net_2273;
  wire net_2287;
  wire net_2288;
  wire net_2289;
  wire net_2291;
  wire net_2293;
  wire net_2295;
  wire net_2297;
  wire net_2298;
  wire net_2309;
  wire net_2315;
  wire net_2322;
  wire net_2327;
  wire net_2330;
  wire net_2331;
  wire net_2332;
  wire net_2333;
  wire net_2334;
  wire net_2336;
  wire net_2337;
  wire net_2338;
  wire net_2339;
  wire net_2340;
  wire net_2342;
  wire net_2343;
  wire net_2345;
  wire net_2347;
  wire net_2348;
  wire net_2349;
  wire net_2350;
  wire net_2351;
  wire net_2352;
  wire net_2353;
  wire net_2354;
  wire net_2355;
  wire net_2356;
  wire net_2357;
  wire net_2358;
  wire net_2359;
  wire net_2360;
  wire net_2361;
  wire net_2362;
  wire net_2364;
  wire net_2365;
  wire net_2366;
  wire net_2367;
  wire net_2368;
  wire net_2369;
  wire net_2370;
  wire net_2371;
  wire net_2396;
  wire net_2398;
  wire net_2399;
  wire net_2400;
  wire net_2401;
  wire net_2402;
  wire net_2403;
  wire net_2407;
  wire net_2444;
  wire net_2446;
  wire net_2448;
  wire net_2456;
  wire net_2478;
  wire net_2485;
  wire net_2488;
  wire net_2489;
  wire net_2490;
  wire net_2491;
  wire net_2492;
  wire net_2493;
  wire net_2497;
  wire net_2498;
  wire net_2501;
  wire net_2503;
  wire net_2520;
  wire net_2521;
  wire net_2522;
  wire net_2523;
  wire net_2524;
  wire net_2526;
  wire net_2528;
  wire net_2529;
  wire net_2530;
  wire net_2531;
  wire net_2533;
  wire net_2534;
  wire net_2535;
  wire net_2544;
  wire net_2546;
  wire net_2548;
  wire net_2553;
  wire net_2554;
  wire net_2555;
  wire net_2556;
  wire net_2557;
  wire net_2558;
  wire net_2559;
  wire net_2560;
  wire net_2561;
  wire net_2562;
  wire net_2563;
  wire net_2564;
  wire net_2565;
  wire net_2566;
  wire net_2567;
  wire net_2568;
  wire net_2572;
  wire net_2573;
  wire net_2574;
  wire net_2575;
  wire net_2576;
  wire net_2577;
  wire net_2578;
  wire net_2579;
  wire net_2604;
  wire net_2605;
  wire net_2606;
  wire net_2607;
  wire net_2608;
  wire net_2609;
  wire net_2610;
  wire net_2611;
  wire net_2657;
  wire net_2660;
  wire net_2665;
  wire net_2670;
  wire net_2702;
  wire net_2703;
  wire net_2719;
  wire net_2720;
  wire net_2721;
  wire net_2781;
  wire net_2782;
  wire net_2783;
  wire net_2784;
  wire net_2785;
  wire net_2786;
  wire net_2787;
  wire net_2813;
  wire net_2814;
  wire net_2815;
  wire net_2816;
  wire net_2817;
  wire net_2818;
  wire net_2819;
  wire net_2820;
  wire net_2861;
  wire net_2864;
  wire net_2868;
  wire net_2870;
  wire net_2872;
  wire net_2873;
  wire net_2878;
  wire net_2893;
  wire net_2913;
  wire net_2920;
  wire net_2926;
  wire net_3025;
  wire net_3026;
  wire net_3027;
  wire net_3028;
  wire net_3029;
  wire net_3030;
  wire net_3031;
  wire net_3032;
  wire net_3092;
  wire net_3137;
  wire net_3139;
  wire net_3151;
  wire net_3157;
  wire net_3158;
  wire net_3218;
  wire net_3219;
  wire net_3220;
  wire net_3221;
  wire net_3222;
  wire net_3223;
  wire net_3224;
  wire net_3225;
  wire net_3250;
  wire net_3251;
  wire net_3252;
  wire net_3253;
  wire net_3254;
  wire net_3255;
  wire net_3256;
  wire net_3300;
  wire net_3304;
  wire net_3306;
  wire net_3308;
  wire net_3344;
  wire net_3348;
  wire net_3350;
  wire net_3351;
  wire net_3354;
  wire net_3356;
  wire net_3362;
  wire net_3365;
  wire net_3380;
  wire net_3382;
  wire net_3383;
  wire net_3385;
  wire net_3386;
  wire net_3388;
  wire net_3389;
  wire net_3390;
  wire net_3392;
  wire net_3393;
  wire net_3394;
  wire net_3395;
  wire net_3397;
  wire net_3399;
  wire net_3400;
  wire net_3402;
  wire net_3407;
  wire net_3408;
  wire net_3409;
  wire net_3410;
  wire net_3411;
  wire net_3412;
  wire net_3413;
  wire net_3414;
  wire net_3415;
  wire net_3416;
  wire net_3417;
  wire net_3418;
  wire net_3419;
  wire net_3420;
  wire net_3421;
  wire net_3422;
  wire net_3424;
  wire net_3425;
  wire net_3426;
  wire net_3427;
  wire net_3428;
  wire net_3429;
  wire net_3430;
  wire net_3431;
  wire net_3457;
  wire net_3458;
  wire net_3459;
  wire net_3463;
  wire net_3514;
  wire net_3553;
  wire net_3556;
  wire net_3559;
  wire net_3562;
  wire net_3580;
  wire net_3582;
  wire net_3583;
  wire net_3585;
  wire net_3587;
  wire net_3589;
  wire net_3590;
  wire net_3592;
  wire net_3594;
  wire net_3595;
  wire net_3597;
  wire net_3598;
  wire net_3600;
  wire net_3606;
  wire net_3607;
  wire net_3611;
  wire net_3613;
  wire net_3614;
  wire net_3615;
  wire net_3616;
  wire net_3617;
  wire net_3618;
  wire net_3619;
  wire net_3620;
  wire net_3621;
  wire net_3622;
  wire net_3623;
  wire net_3624;
  wire net_3625;
  wire net_3626;
  wire net_3627;
  wire net_3628;
  wire net_3632;
  wire net_3633;
  wire net_3634;
  wire net_3635;
  wire net_3636;
  wire net_3637;
  wire net_3638;
  wire net_3639;
  wire net_3664;
  wire net_3665;
  wire net_3668;
  wire net_3670;
  wire net_3731;
  wire net_3746;
  wire net_3758;
  wire net_3841;
  wire net_3842;
  wire net_3843;
  wire net_3844;
  wire net_3845;
  wire net_3846;
  wire net_3847;
  wire net_3873;
  wire net_3878;
  wire net_3880;
  wire net_3965;
  wire net_3976;
  wire net_4086;
  wire net_4087;
  wire net_4091;
  wire net_4092;
  wire net_4312;
  wire net_4315;
  wire net_4423;
  wire net_4425;
  wire net_4427;
  wire net_4429;
  wire net_4431;
  wire net_4433;
  wire net_4435;
  wire net_4540;
  wire net_4544;
  wire net_4545;
  wire net_4650;
  wire net_4653;
  wire net_4654;
  wire net_4658;
  wire net_4660;
  wire net_4768;
  wire net_4879;
  wire net_4880;
  wire net_4881;
  wire net_4900;
  wire net_4959;
  wire net_4960;
  wire net_4961;
  wire net_4962;
  wire net_4963;
  wire net_4964;
  wire net_4965;
  wire net_4966;
  wire net_5039;
  wire net_5088;
  wire net_5091;
  wire net_5093;
  wire net_5095;
  wire net_5097;
  wire net_5117;
  wire net_5118;
  wire net_5120;
  wire net_5122;
  wire net_5123;
  wire net_5125;
  wire net_5126;
  wire net_5127;
  wire net_5128;
  wire net_5133;
  wire net_5134;
  wire net_5140;
  wire net_5141;
  wire net_5142;
  wire net_5144;
  wire net_5146;
  wire net_5148;
  wire net_5149;
  wire net_5150;
  wire net_5151;
  wire net_5152;
  wire net_5153;
  wire net_5154;
  wire net_5155;
  wire net_5156;
  wire net_5157;
  wire net_5158;
  wire net_5159;
  wire net_5160;
  wire net_5161;
  wire net_5162;
  wire net_5163;
  wire net_5165;
  wire net_5166;
  wire net_5167;
  wire net_5168;
  wire net_5169;
  wire net_5170;
  wire net_5171;
  wire net_5172;
  wire net_5260;
  wire net_5298;
  wire net_5299;
  wire net_5302;
  wire net_5323;
  wire net_5325;
  wire net_5326;
  wire net_5327;
  wire net_5328;
  wire net_5329;
  wire net_5330;
  wire net_5331;
  wire net_5332;
  wire net_5336;
  wire net_5340;
  wire net_5341;
  wire net_5342;
  wire net_5344;
  wire net_5345;
  wire net_5346;
  wire net_5354;
  wire net_5355;
  wire net_5356;
  wire net_5357;
  wire net_5358;
  wire net_5359;
  wire net_5360;
  wire net_5361;
  wire net_5362;
  wire net_5363;
  wire net_5364;
  wire net_5365;
  wire net_5366;
  wire net_5367;
  wire net_5368;
  wire net_5369;
  wire net_5373;
  wire net_5374;
  wire net_5375;
  wire net_5376;
  wire net_5377;
  wire net_5378;
  wire net_5379;
  wire net_5380;
  wire net_5453;
  wire net_5472;
  wire net_5497;
  wire net_5499;
  wire net_5511;
  wire net_5582;
  wire net_5583;
  wire net_5584;
  wire net_5585;
  wire net_5586;
  wire net_5587;
  wire net_5588;
  wire net_5683;
  wire net_6673;
  wire net_6674;
  wire net_6676;
  wire net_6678;
  wire net_6680;
  wire net_6717;
  wire net_6720;
  wire net_6721;
  wire net_6726;
  wire net_6727;
  wire net_6730;
  wire net_6745;
  wire net_6760;
  wire net_6761;
  wire net_6763;
  wire net_6778;
  wire net_6779;
  wire net_6781;
  wire net_6784;
  wire net_6792;
  wire net_6795;
  wire net_6796;
  wire net_6825;
  wire net_6826;
  wire net_6827;
  wire net_6828;
  wire net_6829;
  wire net_6830;
  wire net_6831;
  wire net_6832;
  wire net_6871;
  wire net_6886;
  wire net_6889;
  wire net_6891;
  wire net_6904;
  wire net_6905;
  wire net_6907;
  wire net_6909;
  wire net_6912;
  wire net_6915;
  wire net_6917;
  wire net_6919;
  wire net_6922;
  wire net_6924;
  wire net_6925;
  wire net_6937;
  wire net_6940;
  wire net_6943;
  wire net_6944;
  wire net_6946;
  wire net_6949;
  wire net_6950;
  wire net_6952;
  wire net_6955;
  wire net_6956;
  wire net_6958;
  wire net_6960;
  wire net_6962;
  wire net_6964;
  wire net_6967;
  wire net_6968;
  wire net_6971;
  wire net_6974;
  wire net_6977;
  wire net_6978;
  wire net_6979;
  wire net_6980;
  wire net_6982;
  wire net_6983;
  wire net_7008;
  wire net_7009;
  wire net_7010;
  wire net_7011;
  wire net_7012;
  wire net_7013;
  wire net_7014;
  wire net_7015;
  wire net_7023;
  wire net_7032;
  wire net_7036;
  wire net_7050;
  wire net_7052;
  wire net_7056;
  wire net_7057;
  wire net_7058;
  wire net_7060;
  wire net_7062;
  wire net_7065;
  wire net_7066;
  wire net_7072;
  wire net_7074;
  wire net_7075;
  wire net_7077;
  wire net_7078;
  wire net_7082;
  wire net_7084;
  wire net_7085;
  wire net_7088;
  wire net_7089;
  wire net_7090;
  wire net_7096;
  wire net_7100;
  wire net_7108;
  wire net_7114;
  wire net_7118;
  wire net_7119;
  wire net_7120;
  wire net_7121;
  wire net_7124;
  wire net_7126;
  wire net_7127;
  wire net_7129;
  wire net_7130;
  wire net_7155;
  wire net_7156;
  wire net_7157;
  wire net_7158;
  wire net_7159;
  wire net_7160;
  wire net_7161;
  wire net_7162;
  wire net_7169;
  wire net_7176;
  wire net_7177;
  wire net_7179;
  wire net_7196;
  wire net_7199;
  wire net_7201;
  wire net_7205;
  wire net_7207;
  wire net_7209;
  wire net_7213;
  wire net_7214;
  wire net_7218;
  wire net_7222;
  wire net_7226;
  wire net_7231;
  wire net_7234;
  wire net_7236;
  wire net_7238;
  wire net_7240;
  wire net_7242;
  wire net_7244;
  wire net_7246;
  wire net_7248;
  wire net_7250;
  wire net_7252;
  wire net_7254;
  wire net_7256;
  wire net_7258;
  wire net_7261;
  wire net_7262;
  wire net_7265;
  wire net_7268;
  wire net_7271;
  wire net_7272;
  wire net_7273;
  wire net_7274;
  wire net_7276;
  wire net_7277;
  wire net_7302;
  wire net_7304;
  wire net_7305;
  wire net_7306;
  wire net_7308;
  wire net_7309;
  wire net_7335;
  wire net_7343;
  wire net_7346;
  wire net_7349;
  wire net_7353;
  wire net_7357;
  wire net_7359;
  wire net_7361;
  wire net_7363;
  wire net_7364;
  wire net_7366;
  wire net_7377;
  wire net_7384;
  wire net_7390;
  wire net_7395;
  wire net_7402;
  wire net_7407;
  wire net_7408;
  wire net_7409;
  wire net_7415;
  wire net_7418;
  wire net_7423;
  wire net_7424;
  wire net_7449;
  wire net_7450;
  wire net_7451;
  wire net_7452;
  wire net_7453;
  wire net_7454;
  wire net_7455;
  wire net_7459;
  wire net_7463;
  wire net_7465;
  wire net_7469;
  wire net_7471;
  wire net_7491;
  wire net_7506;
  wire net_7509;
  wire net_7510;
  wire net_7519;
  wire net_7529;
  wire net_7543;
  wire net_7549;
  wire net_7554;
  wire net_7561;
  wire net_7570;
  wire net_7571;
  wire net_7596;
  wire net_7597;
  wire net_7599;
  wire net_7600;
  wire net_7602;
  wire net_7603;
  wire net_7619;
  wire net_7648;
  wire net_7651;
  wire net_7676;
  wire net_7716;
  wire net_7717;
  wire net_7743;
  wire net_7744;
  wire net_7745;
  wire net_7746;
  wire net_7747;
  wire net_7748;
  wire net_7749;
  wire net_7750;
  wire net_7759;
  wire net_7767;
  wire net_7771;
  wire net_7792;
  wire net_7798;
  wire net_7801;
  wire net_7802;
  wire net_7806;
  wire net_7808;
  wire net_7812;
  wire net_7815;
  wire net_7817;
  wire net_7823;
  wire net_7832;
  wire net_7835;
  wire net_7842;
  wire net_7850;
  wire net_7853;
  wire net_7861;
  wire net_7864;
  wire net_7865;
  wire net_7890;
  wire net_7891;
  wire net_7892;
  wire net_7893;
  wire net_7894;
  wire net_7895;
  wire net_7896;
  wire net_7897;
  wire net_7898;
  wire net_7904;
  wire net_7915;
  wire net_7918;
  wire net_7920;
  wire net_7923;
  wire net_7931;
  wire net_7936;
  wire net_7944;
  wire net_7946;
  wire net_7956;
  wire net_7960;
  wire net_7961;
  wire net_7962;
  wire net_7966;
  wire net_7973;
  wire net_7977;
  wire net_7982;
  wire net_7988;
  wire net_7997;
  wire net_8000;
  wire net_8007;
  wire net_8011;
  wire net_8012;
  wire net_8037;
  wire net_8039;
  wire net_8041;
  wire net_8042;
  wire net_8043;
  wire net_8044;
  wire net_8050;
  wire net_8052;
  wire net_8065;
  wire net_8066;
  wire net_8070;
  wire net_8071;
  wire net_8072;
  wire net_8081;
  wire net_8083;
  wire net_8085;
  wire net_8089;
  wire net_8095;
  wire net_8098;
  wire net_8104;
  wire net_8108;
  wire net_8114;
  wire net_8120;
  wire net_8124;
  wire net_8131;
  wire net_8136;
  wire net_8143;
  wire net_8149;
  wire net_8155;
  wire net_8158;
  wire net_8159;
  wire net_8185;
  wire net_8186;
  wire net_8187;
  wire net_8188;
  wire net_8189;
  wire net_8190;
  wire net_8191;
  wire net_8202;
  wire net_8219;
  wire net_8228;
  wire net_8232;
  wire net_8235;
  wire net_8246;
  wire net_8247;
  wire net_8248;
  wire net_8252;
  wire net_8254;
  wire net_8261;
  wire net_8266;
  wire net_8271;
  wire net_8276;
  wire net_8283;
  wire net_8291;
  wire net_8294;
  wire net_8303;
  wire net_8305;
  wire net_8306;
  wire net_8331;
  wire net_8332;
  wire net_8333;
  wire net_8334;
  wire net_8335;
  wire net_8336;
  wire net_8337;
  wire net_8338;
  wire net_8351;
  wire net_8354;
  wire net_8355;
  wire net_8361;
  wire net_8362;
  wire net_8363;
  wire net_8364;
  wire net_8375;
  wire net_8377;
  wire net_8378;
  wire net_8380;
  wire net_8383;
  wire net_8384;
  wire net_8392;
  wire net_8406;
  wire net_8418;
  wire net_8424;
  wire net_8430;
  wire net_8438;
  wire net_8444;
  wire net_8450;
  wire net_8452;
  wire net_8453;
  wire net_8478;
  wire net_8479;
  wire net_8480;
  wire net_8481;
  wire net_8482;
  wire net_8483;
  wire net_8484;
  wire net_8485;
  wire net_8505;
  wire net_8519;
  wire net_8522;
  wire net_8525;
  wire net_8527;
  wire net_8529;
  wire net_8531;
  wire net_8533;
  wire net_8535;
  wire net_8553;
  wire net_8560;
  wire net_8564;
  wire net_8573;
  wire net_8576;
  wire net_8582;
  wire net_8591;
  wire net_8594;
  wire net_8599;
  wire net_8600;
  wire net_8626;
  wire net_8627;
  wire net_8628;
  wire net_8629;
  wire net_8630;
  wire net_8631;
  wire net_8632;
  wire net_8637;
  wire net_8641;
  wire net_8643;
  wire net_8647;
  wire net_8669;
  wire net_8670;
  wire net_8671;
  wire net_8673;
  wire net_8680;
  wire net_8683;
  wire net_8684;
  wire net_8689;
  wire net_8700;
  wire net_8707;
  wire net_8714;
  wire net_8719;
  wire net_8726;
  wire net_8730;
  wire net_8735;
  wire net_8743;
  wire net_8746;
  wire net_8747;
  wire net_8773;
  wire net_8774;
  wire net_8775;
  wire net_8776;
  wire net_8777;
  wire net_8778;
  wire net_8779;
  wire net_8785;
  wire net_8802;
  wire net_8813;
  wire net_8824;
  wire net_8827;
  wire net_8829;
  wire net_8830;
  wire net_8835;
  wire net_8838;
  wire net_8841;
  wire net_8846;
  wire net_8854;
  wire net_8861;
  wire net_8866;
  wire net_8870;
  wire net_8879;
  wire net_8882;
  wire net_8891;
  wire net_8893;
  wire net_8894;
  wire net_8919;
  wire net_8920;
  wire net_8921;
  wire net_8922;
  wire net_8923;
  wire net_8924;
  wire net_8925;
  wire net_8926;
  wire net_8936;
  wire net_8965;
  wire net_8977;
  wire net_8981;
  wire net_8982;
  wire net_8984;
  wire net_8988;
  wire net_8989;
  wire net_8996;
  wire net_9001;
  wire net_9008;
  wire net_9014;
  wire net_9018;
  wire net_9024;
  wire net_9030;
  wire net_9040;
  wire net_9041;
  wire net_9068;
  wire net_9071;
  wire net_9073;
  wire net_9082;
  wire net_9097;
  wire net_9107;
  wire net_9108;
  wire net_9111;
  wire net_9130;
  wire net_9146;
  wire net_9154;
  wire net_9159;
  wire net_9182;
  wire net_9187;
  wire net_9188;
  wire net_9213;
  wire net_9214;
  wire net_9217;
  wire net_9219;
  wire net_9220;
  wire net_9256;
  wire net_9261;
  wire net_9267;
  wire net_9281;
  wire net_9289;
  wire net_9295;
  wire net_9311;
  wire net_9323;
  wire net_9334;
  wire net_9335;
  wire net_9360;
  wire net_9361;
  wire net_9363;
  wire net_9364;
  wire net_9365;
  wire net_9366;
  wire net_9367;
  wire net_9387;
  wire net_9402;
  wire net_9407;
  wire net_9416;
  wire net_9436;
  wire net_9465;
  wire net_9476;
  wire net_9481;
  wire net_9482;
  wire net_9508;
  wire net_9510;
  wire net_9511;
  wire net_9512;
  wire net_9514;
  wire net_9554;
  wire net_9560;
  wire net_9564;
  wire net_9576;
  wire net_9590;
  wire net_9596;
  wire net_9617;
  wire net_9625;
  wire net_9628;
  wire net_9629;
  wire net_9655;
  wire net_9658;
  wire net_9700;
  wire net_9721;
  wire net_9729;
  wire net_9748;
  wire net_9775;
  wire net_9776;
  wire net_9801;
  wire net_9806;
  wire net_9843;
  wire net_9848;
  wire net_9851;
  wire net_9882;
  wire net_9905;
  wire net_9913;
  wire net_9922;
  wire net_9923;
  wire net_9952;
  wire net_10015;
  wire net_10037;
  wire net_10069;
  wire net_10070;
  wire net_11229;
  wire net_11230;
  wire net_11231;
  wire net_11232;
  wire net_11235;
  wire net_11236;
  wire net_11272;
  wire net_11278;
  wire net_11279;
  wire net_11283;
  wire net_11293;
  wire net_11294;
  wire net_11295;
  wire net_11302;
  wire net_11304;
  wire net_11305;
  wire net_11307;
  wire net_11310;
  wire net_11322;
  wire net_11323;
  wire net_11324;
  wire net_11325;
  wire net_11336;
  wire net_11346;
  wire net_11348;
  wire net_11351;
  wire net_11352;
  wire net_11357;
  wire net_11358;
  wire net_11359;
  wire net_11360;
  wire net_11361;
  wire net_11362;
  wire net_11363;
  wire net_11364;
  wire net_11370;
  wire net_11374;
  wire net_11378;
  wire net_11380;
  wire net_11417;
  wire net_11421;
  wire net_11423;
  wire net_11435;
  wire net_11436;
  wire net_11437;
  wire net_11438;
  wire net_11439;
  wire net_11440;
  wire net_11442;
  wire net_11444;
  wire net_11445;
  wire net_11446;
  wire net_11447;
  wire net_11448;
  wire net_11449;
  wire net_11451;
  wire net_11452;
  wire net_11454;
  wire net_11455;
  wire net_11462;
  wire net_11465;
  wire net_11469;
  wire net_11474;
  wire net_11475;
  wire net_11476;
  wire net_11479;
  wire net_11480;
  wire net_11481;
  wire net_11482;
  wire net_11485;
  wire net_11486;
  wire net_11487;
  wire net_11488;
  wire net_11492;
  wire net_11497;
  wire net_11498;
  wire net_11499;
  wire net_11500;
  wire net_11503;
  wire net_11505;
  wire net_11506;
  wire net_11509;
  wire net_11510;
  wire net_11511;
  wire net_11514;
  wire net_11515;
  wire net_11516;
  wire net_11517;
  wire net_11518;
  wire net_11519;
  wire net_11520;
  wire net_11521;
  wire net_11522;
  wire net_11523;
  wire net_11528;
  wire net_11536;
  wire net_11538;
  wire net_11541;
  wire net_11543;
  wire net_11548;
  wire net_11558;
  wire net_11560;
  wire net_11561;
  wire net_11562;
  wire net_11563;
  wire net_11564;
  wire net_11565;
  wire net_11567;
  wire net_11569;
  wire net_11570;
  wire net_11572;
  wire net_11573;
  wire net_11575;
  wire net_11585;
  wire net_11586;
  wire net_11588;
  wire net_11590;
  wire net_11591;
  wire net_11593;
  wire net_11596;
  wire net_11597;
  wire net_11598;
  wire net_11603;
  wire net_11611;
  wire net_11614;
  wire net_11615;
  wire net_11616;
  wire net_11620;
  wire net_11621;
  wire net_11622;
  wire net_11623;
  wire net_11626;
  wire net_11627;
  wire net_11628;
  wire net_11629;
  wire net_11632;
  wire net_11633;
  wire net_11634;
  wire net_11635;
  wire net_11637;
  wire net_11638;
  wire net_11639;
  wire net_11641;
  wire net_11642;
  wire net_11643;
  wire net_11644;
  wire net_11645;
  wire net_11646;
  wire net_11667;
  wire net_11668;
  wire net_11672;
  wire net_11680;
  wire net_11682;
  wire net_11683;
  wire net_11684;
  wire net_11686;
  wire net_11690;
  wire net_11692;
  wire net_11693;
  wire net_11695;
  wire net_11696;
  wire net_11699;
  wire net_11702;
  wire net_11704;
  wire net_11706;
  wire net_11707;
  wire net_11708;
  wire net_11709;
  wire net_11710;
  wire net_11713;
  wire net_11714;
  wire net_11715;
  wire net_11716;
  wire net_11719;
  wire net_11720;
  wire net_11722;
  wire net_11728;
  wire net_11731;
  wire net_11732;
  wire net_11733;
  wire net_11734;
  wire net_11737;
  wire net_11738;
  wire net_11739;
  wire net_11740;
  wire net_11745;
  wire net_11749;
  wire net_11750;
  wire net_11751;
  wire net_11755;
  wire net_11756;
  wire net_11758;
  wire net_11760;
  wire net_11761;
  wire net_11762;
  wire net_11763;
  wire net_11764;
  wire net_11766;
  wire net_11767;
  wire net_11768;
  wire net_11769;
  wire net_11775;
  wire net_11776;
  wire net_11778;
  wire net_11787;
  wire net_11788;
  wire net_11790;
  wire net_11795;
  wire net_11796;
  wire net_11809;
  wire net_11816;
  wire net_11819;
  wire net_11821;
  wire net_11825;
  wire net_11829;
  wire net_11831;
  wire net_11833;
  wire net_11838;
  wire net_11848;
  wire net_11850;
  wire net_11851;
  wire net_11855;
  wire net_11862;
  wire net_11875;
  wire net_11878;
  wire net_11883;
  wire net_11884;
  wire net_11885;
  wire net_11886;
  wire net_11888;
  wire net_11889;
  wire net_11890;
  wire net_11891;
  wire net_11892;
  wire net_11898;
  wire net_11902;
  wire net_11903;
  wire net_11904;
  wire net_11912;
  wire net_11917;
  wire net_11919;
  wire net_11930;
  wire net_11941;
  wire net_11943;
  wire net_11950;
  wire net_11954;
  wire net_11956;
  wire net_11957;
  wire net_11962;
  wire net_11967;
  wire net_11973;
  wire net_11979;
  wire net_11983;
  wire net_11991;
  wire net_11995;
  wire net_12006;
  wire net_12007;
  wire net_12009;
  wire net_12010;
  wire net_12011;
  wire net_12012;
  wire net_12013;
  wire net_12014;
  wire net_12015;
  wire net_12021;
  wire net_12022;
  wire net_12050;
  wire net_12053;
  wire net_12054;
  wire net_12056;
  wire net_12065;
  wire net_12067;
  wire net_12071;
  wire net_12073;
  wire net_12077;
  wire net_12083;
  wire net_12088;
  wire net_12089;
  wire net_12090;
  wire net_12091;
  wire net_12100;
  wire net_12106;
  wire net_12120;
  wire net_12124;
  wire net_12128;
  wire net_12129;
  wire net_12131;
  wire net_12133;
  wire net_12135;
  wire net_12138;
  wire net_12156;
  wire net_12160;
  wire net_12163;
  wire net_12164;
  wire net_12165;
  wire net_12166;
  wire net_12172;
  wire net_12174;
  wire net_12175;
  wire net_12176;
  wire net_12177;
  wire net_12178;
  wire net_12179;
  wire net_12180;
  wire net_12181;
  wire net_12182;
  wire net_12183;
  wire net_12184;
  wire net_12186;
  wire net_12187;
  wire net_12190;
  wire net_12193;
  wire net_12194;
  wire net_12201;
  wire net_12205;
  wire net_12206;
  wire net_12207;
  wire net_12208;
  wire net_12211;
  wire net_12212;
  wire net_12213;
  wire net_12214;
  wire net_12220;
  wire net_12223;
  wire net_12224;
  wire net_12225;
  wire net_12226;
  wire net_12229;
  wire net_12230;
  wire net_12231;
  wire net_12232;
  wire net_12238;
  wire net_12241;
  wire net_12249;
  wire net_12251;
  wire net_12252;
  wire net_12255;
  wire net_12256;
  wire net_12257;
  wire net_12258;
  wire net_12259;
  wire net_12260;
  wire net_12261;
  wire net_12274;
  wire net_12276;
  wire net_12277;
  wire net_12284;
  wire net_12288;
  wire net_12295;
  wire net_12297;
  wire net_12299;
  wire net_12300;
  wire net_12302;
  wire net_12308;
  wire net_12312;
  wire net_12319;
  wire net_12328;
  wire net_12334;
  wire net_12343;
  wire net_12346;
  wire net_12352;
  wire net_12358;
  wire net_12364;
  wire net_12373;
  wire net_12375;
  wire net_12376;
  wire net_12377;
  wire net_12378;
  wire net_12379;
  wire net_12380;
  wire net_12381;
  wire net_12382;
  wire net_12383;
  wire net_12384;
  wire net_12389;
  wire net_12399;
  wire net_12404;
  wire net_12407;
  wire net_12411;
  wire net_12419;
  wire net_12432;
  wire net_12433;
  wire net_12436;
  wire net_12439;
  wire net_12442;
  wire net_12443;
  wire net_12446;
  wire net_12452;
  wire net_12464;
  wire net_12475;
  wire net_12476;
  wire net_12477;
  wire net_12483;
  wire net_12488;
  wire net_12496;
  wire net_12497;
  wire net_12498;
  wire net_12500;
  wire net_12501;
  wire net_12502;
  wire net_12503;
  wire net_12504;
  wire net_12505;
  wire net_12506;
  wire net_12507;
  wire net_12516;
  wire net_12525;
  wire net_12530;
  wire net_12534;
  wire net_12541;
  wire net_12542;
  wire net_12544;
  wire net_12546;
  wire net_12553;
  wire net_12554;
  wire net_12556;
  wire net_12559;
  wire net_12563;
  wire net_12564;
  wire net_12565;
  wire net_12566;
  wire net_12567;
  wire net_12568;
  wire net_12569;
  wire net_12570;
  wire net_12573;
  wire net_12575;
  wire net_12576;
  wire net_12579;
  wire net_12581;
  wire net_12582;
  wire net_12583;
  wire net_12585;
  wire net_12587;
  wire net_12588;
  wire net_12589;
  wire net_12591;
  wire net_12593;
  wire net_12594;
  wire net_12595;
  wire net_12597;
  wire net_12599;
  wire net_12600;
  wire net_12601;
  wire net_12603;
  wire net_12605;
  wire net_12606;
  wire net_12607;
  wire net_12609;
  wire net_12611;
  wire net_12612;
  wire net_12613;
  wire net_12615;
  wire net_12617;
  wire net_12618;
  wire net_12619;
  wire net_12621;
  wire net_12622;
  wire net_12624;
  wire net_12625;
  wire net_12626;
  wire net_12627;
  wire net_12628;
  wire net_12629;
  wire net_12630;
  wire net_12653;
  wire net_12654;
  wire net_12658;
  wire net_12659;
  wire net_12667;
  wire net_12669;
  wire net_12681;
  wire net_12683;
  wire net_12685;
  wire net_12688;
  wire net_12690;
  wire net_12692;
  wire net_12695;
  wire net_12696;
  wire net_12698;
  wire net_12699;
  wire net_12700;
  wire net_12702;
  wire net_12704;
  wire net_12705;
  wire net_12706;
  wire net_12708;
  wire net_12710;
  wire net_12711;
  wire net_12712;
  wire net_12714;
  wire net_12716;
  wire net_12717;
  wire net_12718;
  wire net_12720;
  wire net_12722;
  wire net_12723;
  wire net_12724;
  wire net_12726;
  wire net_12728;
  wire net_12729;
  wire net_12730;
  wire net_12732;
  wire net_12734;
  wire net_12735;
  wire net_12736;
  wire net_12738;
  wire net_12740;
  wire net_12741;
  wire net_12742;
  wire net_12744;
  wire net_12745;
  wire net_12747;
  wire net_12748;
  wire net_12749;
  wire net_12750;
  wire net_12751;
  wire net_12752;
  wire net_12753;
  wire net_12758;
  wire net_12761;
  wire net_12770;
  wire net_12775;
  wire net_12779;
  wire net_12781;
  wire net_12782;
  wire net_12790;
  wire net_12793;
  wire net_12798;
  wire net_12802;
  wire net_12804;
  wire net_12810;
  wire net_12812;
  wire net_12814;
  wire net_12816;
  wire net_12818;
  wire net_12820;
  wire net_12822;
  wire net_12823;
  wire net_12828;
  wire net_12832;
  wire net_12840;
  wire net_12844;
  wire net_12853;
  wire net_12857;
  wire net_12863;
  wire net_12865;
  wire net_12867;
  wire net_12868;
  wire net_12869;
  wire net_12870;
  wire net_12871;
  wire net_12872;
  wire net_12873;
  wire net_12874;
  wire net_12875;
  wire net_12876;
  wire net_12882;
  wire net_12883;
  wire net_12884;
  wire net_12887;
  wire net_12889;
  wire net_12892;
  wire net_12894;
  wire net_12895;
  wire net_12898;
  wire net_12899;
  wire net_12900;
  wire net_12903;
  wire net_12913;
  wire net_12919;
  wire net_12920;
  wire net_12925;
  wire net_12927;
  wire net_12928;
  wire net_12931;
  wire net_12932;
  wire net_12934;
  wire net_12935;
  wire net_12942;
  wire net_12944;
  wire net_12945;
  wire net_12948;
  wire net_12950;
  wire net_12951;
  wire net_12952;
  wire net_12956;
  wire net_12957;
  wire net_12958;
  wire net_12962;
  wire net_12967;
  wire net_12975;
  wire net_12979;
  wire net_12982;
  wire net_12985;
  wire net_12990;
  wire net_12991;
  wire net_12993;
  wire net_12994;
  wire net_12995;
  wire net_12996;
  wire net_12997;
  wire net_12998;
  wire net_12999;
  wire net_13006;
  wire net_13016;
  wire net_13017;
  wire net_13034;
  wire net_13035;
  wire net_13036;
  wire net_13037;
  wire net_13039;
  wire net_13040;
  wire net_13043;
  wire net_13055;
  wire net_13060;
  wire net_13062;
  wire net_13063;
  wire net_13065;
  wire net_13067;
  wire net_13068;
  wire net_13071;
  wire net_13073;
  wire net_13074;
  wire net_13075;
  wire net_13079;
  wire net_13080;
  wire net_13081;
  wire net_13084;
  wire net_13085;
  wire net_13086;
  wire net_13090;
  wire net_13097;
  wire net_13105;
  wire net_13111;
  wire net_13113;
  wire net_13114;
  wire net_13115;
  wire net_13116;
  wire net_13117;
  wire net_13118;
  wire net_13119;
  wire net_13120;
  wire net_13121;
  wire net_13122;
  wire net_13129;
  wire net_13141;
  wire net_13148;
  wire net_13158;
  wire net_13163;
  wire net_13164;
  wire net_13166;
  wire net_13173;
  wire net_13174;
  wire net_13183;
  wire net_13187;
  wire net_13189;
  wire net_13198;
  wire net_13203;
  wire net_13207;
  wire net_13214;
  wire net_13219;
  wire net_13227;
  wire net_13233;
  wire net_13236;
  wire net_13237;
  wire net_13238;
  wire net_13240;
  wire net_13241;
  wire net_13242;
  wire net_13243;
  wire net_13244;
  wire net_13245;
  wire net_13264;
  wire net_13291;
  wire net_13294;
  wire net_13301;
  wire net_13324;
  wire net_13345;
  wire net_13356;
  wire net_13359;
  wire net_13360;
  wire net_13361;
  wire net_13365;
  wire net_13366;
  wire net_13367;
  wire net_13368;
  wire net_13388;
  wire net_13403;
  wire net_13407;
  wire net_13408;
  wire net_13409;
  wire net_13421;
  wire net_13436;
  wire net_13444;
  wire net_13460;
  wire net_13472;
  wire net_13479;
  wire net_13482;
  wire net_13483;
  wire net_13486;
  wire net_13489;
  wire net_13519;
  wire net_13528;
  wire net_13529;
  wire net_13531;
  wire net_13533;
  wire net_13537;
  wire net_13538;
  wire net_13540;
  wire net_13560;
  wire net_13567;
  wire net_13576;
  wire net_13583;
  wire net_13591;
  wire net_13596;
  wire net_13600;
  wire net_13605;
  wire net_13606;
  wire net_13608;
  wire net_13631;
  wire net_13650;
  wire net_13652;
  wire net_13653;
  wire net_13655;
  wire net_13672;
  wire net_13690;
  wire net_13700;
  wire net_13708;
  wire net_13711;
  wire net_13723;
  wire net_13728;
  wire net_13729;
  wire net_13735;
  wire net_13736;
  wire net_13776;
  wire net_13779;
  wire net_13810;
  wire net_13829;
  wire net_13851;
  wire net_13852;
  wire net_13856;
  wire net_13897;
  wire net_13920;
  wire net_13928;
  wire net_13959;
  wire net_13974;
  wire net_13975;
  wire net_14026;
  wire net_14074;
  wire net_14097;
  wire net_14098;
  wire net_15060;
  wire net_15062;
  wire net_15063;
  wire net_15064;
  wire net_15065;
  wire net_15066;
  wire net_15067;
  wire net_15103;
  wire net_15104;
  wire net_15106;
  wire net_15110;
  wire net_15115;
  wire net_15118;
  wire net_15119;
  wire net_15120;
  wire net_15121;
  wire net_15122;
  wire net_15124;
  wire net_15126;
  wire net_15127;
  wire net_15129;
  wire net_15131;
  wire net_15132;
  wire net_15133;
  wire net_15135;
  wire net_15136;
  wire net_15137;
  wire net_15138;
  wire net_15141;
  wire net_15142;
  wire net_15143;
  wire net_15147;
  wire net_15148;
  wire net_15149;
  wire net_15150;
  wire net_15153;
  wire net_15154;
  wire net_15155;
  wire net_15156;
  wire net_15171;
  wire net_15173;
  wire net_15177;
  wire net_15178;
  wire net_15179;
  wire net_15180;
  wire net_15181;
  wire net_15182;
  wire net_15183;
  wire net_15189;
  wire net_15190;
  wire net_15191;
  wire net_15192;
  wire net_15193;
  wire net_15194;
  wire net_15195;
  wire net_15208;
  wire net_15229;
  wire net_15234;
  wire net_15242;
  wire net_15243;
  wire net_15244;
  wire net_15247;
  wire net_15249;
  wire net_15250;
  wire net_15265;
  wire net_15268;
  wire net_15269;
  wire net_15270;
  wire net_15273;
  wire net_15274;
  wire net_15279;
  wire net_15280;
  wire net_15282;
  wire net_15283;
  wire net_15284;
  wire net_15285;
  wire net_15286;
  wire net_15289;
  wire net_15290;
  wire net_15291;
  wire net_15292;
  wire net_15293;
  wire net_15294;
  wire net_15295;
  wire net_15296;
  wire net_15298;
  wire net_15299;
  wire net_15300;
  wire net_15301;
  wire net_15304;
  wire net_15305;
  wire net_15306;
  wire net_15307;
  wire net_15311;
  wire net_15312;
  wire net_15313;
  wire net_15316;
  wire net_15317;
  wire net_15318;
  wire net_15319;
  wire net_15322;
  wire net_15323;
  wire net_15325;
  wire net_15328;
  wire net_15329;
  wire net_15330;
  wire net_15331;
  wire net_15335;
  wire net_15337;
  wire net_15341;
  wire net_15342;
  wire net_15343;
  wire net_15344;
  wire net_15345;
  wire net_15346;
  wire net_15347;
  wire net_15348;
  wire net_15349;
  wire net_15350;
  wire net_15351;
  wire net_15352;
  wire net_15353;
  wire net_15354;
  wire net_15365;
  wire net_15369;
  wire net_15390;
  wire net_15391;
  wire net_15392;
  wire net_15394;
  wire net_15395;
  wire net_15397;
  wire net_15398;
  wire net_15399;
  wire net_15400;
  wire net_15402;
  wire net_15404;
  wire net_15406;
  wire net_15407;
  wire net_15408;
  wire net_15409;
  wire net_15410;
  wire net_15412;
  wire net_15414;
  wire net_15415;
  wire net_15416;
  wire net_15417;
  wire net_15421;
  wire net_15422;
  wire net_15423;
  wire net_15424;
  wire net_15427;
  wire net_15428;
  wire net_15429;
  wire net_15430;
  wire net_15433;
  wire net_15434;
  wire net_15439;
  wire net_15440;
  wire net_15441;
  wire net_15442;
  wire net_15445;
  wire net_15447;
  wire net_15448;
  wire net_15451;
  wire net_15452;
  wire net_15453;
  wire net_15454;
  wire net_15457;
  wire net_15458;
  wire net_15459;
  wire net_15460;
  wire net_15463;
  wire net_15464;
  wire net_15465;
  wire net_15466;
  wire net_15467;
  wire net_15468;
  wire net_15469;
  wire net_15470;
  wire net_15471;
  wire net_15472;
  wire net_15473;
  wire net_15474;
  wire net_15475;
  wire net_15476;
  wire net_15488;
  wire net_15490;
  wire net_15511;
  wire net_15514;
  wire net_15516;
  wire net_15518;
  wire net_15519;
  wire net_15522;
  wire net_15523;
  wire net_15524;
  wire net_15525;
  wire net_15526;
  wire net_15527;
  wire net_15530;
  wire net_15533;
  wire net_15536;
  wire net_15544;
  wire net_15545;
  wire net_15546;
  wire net_15547;
  wire net_15556;
  wire net_15557;
  wire net_15564;
  wire net_15568;
  wire net_15569;
  wire net_15570;
  wire net_15574;
  wire net_15575;
  wire net_15577;
  wire net_15583;
  wire net_15587;
  wire net_15589;
  wire net_15591;
  wire net_15592;
  wire net_15593;
  wire net_15594;
  wire net_15595;
  wire net_15596;
  wire net_15597;
  wire net_15598;
  wire net_15599;
  wire net_15600;
  wire net_15606;
  wire net_15608;
  wire net_15622;
  wire net_15625;
  wire net_15638;
  wire net_15640;
  wire net_15642;
  wire net_15644;
  wire net_15648;
  wire net_15651;
  wire net_15653;
  wire net_15655;
  wire net_15660;
  wire net_15668;
  wire net_15670;
  wire net_15674;
  wire net_15682;
  wire net_15692;
  wire net_15694;
  wire net_15697;
  wire net_15705;
  wire net_15709;
  wire net_15714;
  wire net_15715;
  wire net_15716;
  wire net_15717;
  wire net_15718;
  wire net_15719;
  wire net_15720;
  wire net_15721;
  wire net_15722;
  wire net_15723;
  wire net_15729;
  wire net_15730;
  wire net_15737;
  wire net_15739;
  wire net_15746;
  wire net_15748;
  wire net_15761;
  wire net_15762;
  wire net_15765;
  wire net_15766;
  wire net_15767;
  wire net_15770;
  wire net_15772;
  wire net_15774;
  wire net_15775;
  wire net_15776;
  wire net_15781;
  wire net_15783;
  wire net_15784;
  wire net_15791;
  wire net_15797;
  wire net_15808;
  wire net_15814;
  wire net_15815;
  wire net_15816;
  wire net_15817;
  wire net_15820;
  wire net_15827;
  wire net_15828;
  wire net_15829;
  wire net_15835;
  wire net_15836;
  wire net_15837;
  wire net_15839;
  wire net_15840;
  wire net_15841;
  wire net_15842;
  wire net_15843;
  wire net_15844;
  wire net_15845;
  wire net_15846;
  wire net_15859;
  wire net_15861;
  wire net_15882;
  wire net_15883;
  wire net_15884;
  wire net_15885;
  wire net_15886;
  wire net_15888;
  wire net_15889;
  wire net_15890;
  wire net_15891;
  wire net_15892;
  wire net_15894;
  wire net_15895;
  wire net_15912;
  wire net_15914;
  wire net_15915;
  wire net_15918;
  wire net_15920;
  wire net_15921;
  wire net_15922;
  wire net_15924;
  wire net_15926;
  wire net_15927;
  wire net_15928;
  wire net_15930;
  wire net_15932;
  wire net_15933;
  wire net_15934;
  wire net_15936;
  wire net_15938;
  wire net_15939;
  wire net_15940;
  wire net_15942;
  wire net_15944;
  wire net_15945;
  wire net_15946;
  wire net_15952;
  wire net_15956;
  wire net_15957;
  wire net_15960;
  wire net_15961;
  wire net_15969;
  wire net_16003;
  wire net_16005;
  wire net_16013;
  wire net_16020;
  wire net_16023;
  wire net_16029;
  wire net_16038;
  wire net_16051;
  wire net_16060;
  wire net_16061;
  wire net_16063;
  wire net_16079;
  wire net_16082;
  wire net_16083;
  wire net_16085;
  wire net_16086;
  wire net_16087;
  wire net_16088;
  wire net_16089;
  wire net_16090;
  wire net_16091;
  wire net_16092;
  wire net_16109;
  wire net_16111;
  wire net_16115;
  wire net_16116;
  wire net_16118;
  wire net_16127;
  wire net_16129;
  wire net_16130;
  wire net_16132;
  wire net_16133;
  wire net_16134;
  wire net_16135;
  wire net_16138;
  wire net_16139;
  wire net_16141;
  wire net_16142;
  wire net_16149;
  wire net_16153;
  wire net_16156;
  wire net_16158;
  wire net_16160;
  wire net_16161;
  wire net_16164;
  wire net_16166;
  wire net_16167;
  wire net_16168;
  wire net_16170;
  wire net_16172;
  wire net_16173;
  wire net_16174;
  wire net_16176;
  wire net_16178;
  wire net_16179;
  wire net_16180;
  wire net_16182;
  wire net_16184;
  wire net_16185;
  wire net_16186;
  wire net_16188;
  wire net_16190;
  wire net_16191;
  wire net_16192;
  wire net_16194;
  wire net_16196;
  wire net_16197;
  wire net_16198;
  wire net_16204;
  wire net_16208;
  wire net_16209;
  wire net_16210;
  wire net_16211;
  wire net_16212;
  wire net_16213;
  wire net_16214;
  wire net_16215;
  wire net_16223;
  wire net_16225;
  wire net_16227;
  wire net_16231;
  wire net_16233;
  wire net_16236;
  wire net_16237;
  wire net_16241;
  wire net_16242;
  wire net_16243;
  wire net_16253;
  wire net_16254;
  wire net_16260;
  wire net_16261;
  wire net_16268;
  wire net_16273;
  wire net_16276;
  wire net_16278;
  wire net_16283;
  wire net_16291;
  wire net_16296;
  wire net_16300;
  wire net_16309;
  wire net_16315;
  wire net_16320;
  wire net_16326;
  wire net_16329;
  wire net_16330;
  wire net_16331;
  wire net_16332;
  wire net_16333;
  wire net_16334;
  wire net_16335;
  wire net_16336;
  wire net_16337;
  wire net_16338;
  wire net_16346;
  wire net_16349;
  wire net_16354;
  wire net_16357;
  wire net_16359;
  wire net_16360;
  wire net_16362;
  wire net_16363;
  wire net_16364;
  wire net_16366;
  wire net_16375;
  wire net_16383;
  wire net_16385;
  wire net_16386;
  wire net_16387;
  wire net_16388;
  wire net_16390;
  wire net_16394;
  wire net_16406;
  wire net_16414;
  wire net_16419;
  wire net_16425;
  wire net_16431;
  wire net_16436;
  wire net_16443;
  wire net_16450;
  wire net_16452;
  wire net_16453;
  wire net_16454;
  wire net_16455;
  wire net_16456;
  wire net_16457;
  wire net_16458;
  wire net_16459;
  wire net_16461;
  wire net_16469;
  wire net_16471;
  wire net_16476;
  wire net_16477;
  wire net_16478;
  wire net_16481;
  wire net_16487;
  wire net_16498;
  wire net_16499;
  wire net_16500;
  wire net_16504;
  wire net_16507;
  wire net_16508;
  wire net_16510;
  wire net_16513;
  wire net_16514;
  wire net_16515;
  wire net_16517;
  wire net_16518;
  wire net_16523;
  wire net_16525;
  wire net_16527;
  wire net_16529;
  wire net_16530;
  wire net_16533;
  wire net_16535;
  wire net_16536;
  wire net_16537;
  wire net_16539;
  wire net_16541;
  wire net_16542;
  wire net_16543;
  wire net_16545;
  wire net_16547;
  wire net_16548;
  wire net_16549;
  wire net_16551;
  wire net_16553;
  wire net_16554;
  wire net_16555;
  wire net_16557;
  wire net_16559;
  wire net_16560;
  wire net_16561;
  wire net_16563;
  wire net_16565;
  wire net_16566;
  wire net_16567;
  wire net_16573;
  wire net_16584;
  wire net_16591;
  wire net_16595;
  wire net_16598;
  wire net_16599;
  wire net_16603;
  wire net_16604;
  wire net_16607;
  wire net_16611;
  wire net_16623;
  wire net_16625;
  wire net_16633;
  wire net_16634;
  wire net_16636;
  wire net_16637;
  wire net_16638;
  wire net_16639;
  wire net_16640;
  wire net_16642;
  wire net_16643;
  wire net_16644;
  wire net_16645;
  wire net_16646;
  wire net_16647;
  wire net_16648;
  wire net_16650;
  wire net_16652;
  wire net_16653;
  wire net_16656;
  wire net_16658;
  wire net_16659;
  wire net_16660;
  wire net_16662;
  wire net_16664;
  wire net_16665;
  wire net_16666;
  wire net_16668;
  wire net_16670;
  wire net_16671;
  wire net_16672;
  wire net_16674;
  wire net_16676;
  wire net_16677;
  wire net_16678;
  wire net_16680;
  wire net_16682;
  wire net_16683;
  wire net_16684;
  wire net_16686;
  wire net_16688;
  wire net_16689;
  wire net_16690;
  wire net_16692;
  wire net_16694;
  wire net_16695;
  wire net_16696;
  wire net_16698;
  wire net_16699;
  wire net_16700;
  wire net_16701;
  wire net_16703;
  wire net_16704;
  wire net_16705;
  wire net_16706;
  wire net_16707;
  wire net_16714;
  wire net_16716;
  wire net_16717;
  wire net_16722;
  wire net_16725;
  wire net_16731;
  wire net_16736;
  wire net_16742;
  wire net_16748;
  wire net_16756;
  wire net_16757;
  wire net_16758;
  wire net_16761;
  wire net_16762;
  wire net_16765;
  wire net_16767;
  wire net_16768;
  wire net_16770;
  wire net_16773;
  wire net_16775;
  wire net_16776;
  wire net_16777;
  wire net_16780;
  wire net_16782;
  wire net_16783;
  wire net_16787;
  wire net_16794;
  wire net_16799;
  wire net_16804;
  wire net_16805;
  wire net_16807;
  wire net_16812;
  wire net_16817;
  wire net_16821;
  wire net_16822;
  wire net_16823;
  wire net_16824;
  wire net_16825;
  wire net_16826;
  wire net_16827;
  wire net_16828;
  wire net_16829;
  wire net_16830;
  wire net_16864;
  wire net_16866;
  wire net_16867;
  wire net_16868;
  wire net_16869;
  wire net_16873;
  wire net_16878;
  wire net_16883;
  wire net_16884;
  wire net_16886;
  wire net_16890;
  wire net_16892;
  wire net_16893;
  wire net_16894;
  wire net_16896;
  wire net_16898;
  wire net_16899;
  wire net_16902;
  wire net_16904;
  wire net_16905;
  wire net_16906;
  wire net_16908;
  wire net_16910;
  wire net_16911;
  wire net_16912;
  wire net_16914;
  wire net_16916;
  wire net_16917;
  wire net_16918;
  wire net_16920;
  wire net_16922;
  wire net_16923;
  wire net_16924;
  wire net_16926;
  wire net_16928;
  wire net_16929;
  wire net_16930;
  wire net_16932;
  wire net_16934;
  wire net_16935;
  wire net_16936;
  wire net_16942;
  wire net_16946;
  wire net_16947;
  wire net_16950;
  wire net_16951;
  wire net_16952;
  wire net_16953;
  wire net_16970;
  wire net_16977;
  wire net_16980;
  wire net_16989;
  wire net_16990;
  wire net_16992;
  wire net_16998;
  wire net_16999;
  wire net_17001;
  wire net_17004;
  wire net_17016;
  wire net_17023;
  wire net_17029;
  wire net_17033;
  wire net_17041;
  wire net_17045;
  wire net_17051;
  wire net_17057;
  wire net_17062;
  wire net_17067;
  wire net_17068;
  wire net_17069;
  wire net_17070;
  wire net_17072;
  wire net_17073;
  wire net_17074;
  wire net_17075;
  wire net_17076;
  wire net_17094;
  wire net_17097;
  wire net_17114;
  wire net_17115;
  wire net_17121;
  wire net_17126;
  wire net_17127;
  wire net_17132;
  wire net_17133;
  wire net_17143;
  wire net_17158;
  wire net_17164;
  wire net_17169;
  wire net_17173;
  wire net_17179;
  wire net_17185;
  wire net_17190;
  wire net_17191;
  wire net_17195;
  wire net_17205;
  wire net_17206;
  wire net_17218;
  wire net_17220;
  wire net_17233;
  wire net_17234;
  wire net_17237;
  wire net_17238;
  wire net_17241;
  wire net_17242;
  wire net_17243;
  wire net_17244;
  wire net_17245;
  wire net_17246;
  wire net_17248;
  wire net_17249;
  wire net_17253;
  wire net_17259;
  wire net_17266;
  wire net_17267;
  wire net_17268;
  wire net_17269;
  wire net_17291;
  wire net_17296;
  wire net_17297;
  wire net_17298;
  wire net_17299;
  wire net_17302;
  wire net_17303;
  wire net_17304;
  wire net_17305;
  wire net_17309;
  wire net_17312;
  wire net_17313;
  wire net_17314;
  wire net_17315;
  wire net_17321;
  wire net_17322;
  wire net_17327;
  wire net_17364;
  wire net_17373;
  wire net_17402;
  wire net_17421;
  wire net_17436;
  wire net_17437;
  wire net_17442;
  wire net_17443;
  wire net_17450;
  wire net_17504;
  wire net_17521;
  wire net_17559;
  wire net_17560;
  wire net_17585;
  wire net_17613;
  wire net_17620;
  wire net_17666;
  wire net_17671;
  wire net_17682;
  wire net_17683;
  wire net_17690;
  wire net_17745;
  wire net_17777;
  wire net_17805;
  wire net_17806;
  wire net_18791;
  wire net_18894;
  wire net_18898;
  wire net_18923;
  wire net_18935;
  wire net_18936;
  wire net_18940;
  wire net_18942;
  wire net_18943;
  wire net_18944;
  wire net_18945;
  wire net_18946;
  wire net_18948;
  wire net_18949;
  wire net_18951;
  wire net_18952;
  wire net_18954;
  wire net_18960;
  wire net_18963;
  wire net_18966;
  wire net_18967;
  wire net_18968;
  wire net_18969;
  wire net_18978;
  wire net_18980;
  wire net_18984;
  wire net_18985;
  wire net_18990;
  wire net_18991;
  wire net_18992;
  wire net_18993;
  wire net_18996;
  wire net_18997;
  wire net_18998;
  wire net_18999;
  wire net_19002;
  wire net_19003;
  wire net_19004;
  wire net_19005;
  wire net_19008;
  wire net_19009;
  wire net_19010;
  wire net_19011;
  wire net_19012;
  wire net_19013;
  wire net_19014;
  wire net_19020;
  wire net_19024;
  wire net_19069;
  wire net_19076;
  wire net_19079;
  wire net_19080;
  wire net_19081;
  wire net_19098;
  wire net_19100;
  wire net_19102;
  wire net_19103;
  wire net_19107;
  wire net_19108;
  wire net_19109;
  wire net_19110;
  wire net_19113;
  wire net_19114;
  wire net_19117;
  wire net_19118;
  wire net_19119;
  wire net_19122;
  wire net_19123;
  wire net_19124;
  wire net_19126;
  wire net_19127;
  wire net_19128;
  wire net_19130;
  wire net_19131;
  wire net_19134;
  wire net_19135;
  wire net_19136;
  wire net_19137;
  wire net_19138;
  wire net_19140;
  wire net_19142;
  wire net_19143;
  wire net_19144;
  wire net_19146;
  wire net_19148;
  wire net_19149;
  wire net_19150;
  wire net_19152;
  wire net_19153;
  wire net_19154;
  wire net_19155;
  wire net_19156;
  wire net_19158;
  wire net_19159;
  wire net_19160;
  wire net_19161;
  wire net_19162;
  wire net_19164;
  wire net_19165;
  wire net_19166;
  wire net_19167;
  wire net_19168;
  wire net_19170;
  wire net_19172;
  wire net_19173;
  wire net_19174;
  wire net_19180;
  wire net_19182;
  wire net_19183;
  wire net_19185;
  wire net_19209;
  wire net_19214;
  wire net_19219;
  wire net_19221;
  wire net_19222;
  wire net_19223;
  wire net_19224;
  wire net_19225;
  wire net_19230;
  wire net_19231;
  wire net_19232;
  wire net_19233;
  wire net_19234;
  wire net_19236;
  wire net_19237;
  wire net_19239;
  wire net_19240;
  wire net_19241;
  wire net_19242;
  wire net_19245;
  wire net_19247;
  wire net_19250;
  wire net_19251;
  wire net_19252;
  wire net_19253;
  wire net_19254;
  wire net_19255;
  wire net_19257;
  wire net_19259;
  wire net_19260;
  wire net_19261;
  wire net_19263;
  wire net_19265;
  wire net_19266;
  wire net_19267;
  wire net_19269;
  wire net_19271;
  wire net_19272;
  wire net_19273;
  wire net_19276;
  wire net_19277;
  wire net_19279;
  wire net_19282;
  wire net_19283;
  wire net_19284;
  wire net_19285;
  wire net_19289;
  wire net_19290;
  wire net_19291;
  wire net_19294;
  wire net_19295;
  wire net_19296;
  wire net_19297;
  wire net_19298;
  wire net_19299;
  wire net_19300;
  wire net_19301;
  wire net_19302;
  wire net_19303;
  wire net_19304;
  wire net_19305;
  wire net_19306;
  wire net_19307;
  wire net_19308;
  wire net_19326;
  wire net_19334;
  wire net_19336;
  wire net_19346;
  wire net_19348;
  wire net_19350;
  wire net_19352;
  wire net_19353;
  wire net_19354;
  wire net_19356;
  wire net_19360;
  wire net_19361;
  wire net_19362;
  wire net_19365;
  wire net_19371;
  wire net_19373;
  wire net_19376;
  wire net_19377;
  wire net_19378;
  wire net_19384;
  wire net_19390;
  wire net_19393;
  wire net_19394;
  wire net_19395;
  wire net_19396;
  wire net_19399;
  wire net_19401;
  wire net_19402;
  wire net_19408;
  wire net_19411;
  wire net_19412;
  wire net_19413;
  wire net_19414;
  wire net_19422;
  wire net_19423;
  wire net_19425;
  wire net_19426;
  wire net_19427;
  wire net_19428;
  wire net_19429;
  wire net_19430;
  wire net_19431;
  wire net_19440;
  wire net_19441;
  wire net_19442;
  wire net_19445;
  wire net_19448;
  wire net_19450;
  wire net_19456;
  wire net_19470;
  wire net_19471;
  wire net_19473;
  wire net_19474;
  wire net_19478;
  wire net_19479;
  wire net_19481;
  wire net_19483;
  wire net_19485;
  wire net_19488;
  wire net_19492;
  wire net_19493;
  wire net_19494;
  wire net_19495;
  wire net_19496;
  wire net_19498;
  wire net_19500;
  wire net_19505;
  wire net_19513;
  wire net_19516;
  wire net_19519;
  wire net_19523;
  wire net_19524;
  wire net_19525;
  wire net_19529;
  wire net_19530;
  wire net_19531;
  wire net_19534;
  wire net_19535;
  wire net_19536;
  wire net_19537;
  wire net_19541;
  wire net_19545;
  wire net_19546;
  wire net_19548;
  wire net_19549;
  wire net_19550;
  wire net_19551;
  wire net_19552;
  wire net_19553;
  wire net_19554;
  wire net_19561;
  wire net_19574;
  wire net_19588;
  wire net_19590;
  wire net_19591;
  wire net_19592;
  wire net_19595;
  wire net_19596;
  wire net_19599;
  wire net_19602;
  wire net_19603;
  wire net_19604;
  wire net_19612;
  wire net_19615;
  wire net_19623;
  wire net_19627;
  wire net_19629;
  wire net_19633;
  wire net_19636;
  wire net_19641;
  wire net_19642;
  wire net_19645;
  wire net_19646;
  wire net_19647;
  wire net_19648;
  wire net_19651;
  wire net_19653;
  wire net_19659;
  wire net_19660;
  wire net_19664;
  wire net_19667;
  wire net_19668;
  wire net_19671;
  wire net_19672;
  wire net_19673;
  wire net_19675;
  wire net_19689;
  wire net_19693;
  wire net_19699;
  wire net_19712;
  wire net_19715;
  wire net_19718;
  wire net_19720;
  wire net_19721;
  wire net_19724;
  wire net_19725;
  wire net_19726;
  wire net_19729;
  wire net_19731;
  wire net_19732;
  wire net_19734;
  wire net_19735;
  wire net_19736;
  wire net_19737;
  wire net_19738;
  wire net_19740;
  wire net_19742;
  wire net_19744;
  wire net_19745;
  wire net_19746;
  wire net_19747;
  wire net_19753;
  wire net_19756;
  wire net_19757;
  wire net_19758;
  wire net_19759;
  wire net_19762;
  wire net_19763;
  wire net_19764;
  wire net_19765;
  wire net_19768;
  wire net_19769;
  wire net_19770;
  wire net_19771;
  wire net_19775;
  wire net_19780;
  wire net_19788;
  wire net_19790;
  wire net_19791;
  wire net_19793;
  wire net_19794;
  wire net_19795;
  wire net_19796;
  wire net_19797;
  wire net_19798;
  wire net_19799;
  wire net_19800;
  wire net_19805;
  wire net_19811;
  wire net_19814;
  wire net_19838;
  wire net_19848;
  wire net_19852;
  wire net_19854;
  wire net_19856;
  wire net_19859;
  wire net_19861;
  wire net_19863;
  wire net_19865;
  wire net_19868;
  wire net_19869;
  wire net_19874;
  wire net_19875;
  wire net_19880;
  wire net_19881;
  wire net_19886;
  wire net_19887;
  wire net_19892;
  wire net_19893;
  wire net_19898;
  wire net_19899;
  wire net_19902;
  wire net_19904;
  wire net_19905;
  wire net_19908;
  wire net_19910;
  wire net_19911;
  wire net_19912;
  wire net_19914;
  wire net_19915;
  wire net_19916;
  wire net_19917;
  wire net_19918;
  wire net_19919;
  wire net_19920;
  wire net_19921;
  wire net_19922;
  wire net_19923;
  wire net_19925;
  wire net_19933;
  wire net_19939;
  wire net_19942;
  wire net_19944;
  wire net_19945;
  wire net_19948;
  wire net_19950;
  wire net_19951;
  wire net_19952;
  wire net_19960;
  wire net_19972;
  wire net_19989;
  wire net_19991;
  wire net_19992;
  wire net_19993;
  wire net_19995;
  wire net_19997;
  wire net_19998;
  wire net_19999;
  wire net_20001;
  wire net_20003;
  wire net_20004;
  wire net_20005;
  wire net_20007;
  wire net_20009;
  wire net_20010;
  wire net_20011;
  wire net_20013;
  wire net_20015;
  wire net_20016;
  wire net_20017;
  wire net_20019;
  wire net_20021;
  wire net_20022;
  wire net_20023;
  wire net_20025;
  wire net_20027;
  wire net_20028;
  wire net_20029;
  wire net_20031;
  wire net_20033;
  wire net_20034;
  wire net_20035;
  wire net_20037;
  wire net_20038;
  wire net_20039;
  wire net_20040;
  wire net_20041;
  wire net_20042;
  wire net_20043;
  wire net_20044;
  wire net_20045;
  wire net_20046;
  wire net_20054;
  wire net_20058;
  wire net_20062;
  wire net_20063;
  wire net_20065;
  wire net_20066;
  wire net_20067;
  wire net_20069;
  wire net_20070;
  wire net_20071;
  wire net_20073;
  wire net_20075;
  wire net_20101;
  wire net_20111;
  wire net_20112;
  wire net_20114;
  wire net_20115;
  wire net_20116;
  wire net_20118;
  wire net_20120;
  wire net_20121;
  wire net_20122;
  wire net_20124;
  wire net_20126;
  wire net_20127;
  wire net_20128;
  wire net_20130;
  wire net_20132;
  wire net_20133;
  wire net_20134;
  wire net_20136;
  wire net_20138;
  wire net_20139;
  wire net_20140;
  wire net_20142;
  wire net_20144;
  wire net_20145;
  wire net_20146;
  wire net_20148;
  wire net_20150;
  wire net_20151;
  wire net_20152;
  wire net_20155;
  wire net_20156;
  wire net_20158;
  wire net_20160;
  wire net_20161;
  wire net_20162;
  wire net_20163;
  wire net_20164;
  wire net_20165;
  wire net_20166;
  wire net_20167;
  wire net_20168;
  wire net_20169;
  wire net_20181;
  wire net_20186;
  wire net_20187;
  wire net_20189;
  wire net_20190;
  wire net_20191;
  wire net_20195;
  wire net_20197;
  wire net_20204;
  wire net_20205;
  wire net_20207;
  wire net_20213;
  wire net_20215;
  wire net_20220;
  wire net_20228;
  wire net_20232;
  wire net_20237;
  wire net_20242;
  wire net_20251;
  wire net_20255;
  wire net_20262;
  wire net_20266;
  wire net_20274;
  wire net_20281;
  wire net_20283;
  wire net_20284;
  wire net_20285;
  wire net_20286;
  wire net_20287;
  wire net_20288;
  wire net_20289;
  wire net_20290;
  wire net_20291;
  wire net_20292;
  wire net_20306;
  wire net_20309;
  wire net_20311;
  wire net_20312;
  wire net_20313;
  wire net_20316;
  wire net_20317;
  wire net_20319;
  wire net_20333;
  wire net_20337;
  wire net_20341;
  wire net_20344;
  wire net_20348;
  wire net_20350;
  wire net_20352;
  wire net_20362;
  wire net_20367;
  wire net_20371;
  wire net_20380;
  wire net_20383;
  wire net_20391;
  wire net_20404;
  wire net_20405;
  wire net_20406;
  wire net_20408;
  wire net_20409;
  wire net_20410;
  wire net_20411;
  wire net_20412;
  wire net_20413;
  wire net_20414;
  wire net_20415;
  wire net_20422;
  wire net_20423;
  wire net_20426;
  wire net_20429;
  wire net_20435;
  wire net_20437;
  wire net_20443;
  wire net_20449;
  wire net_20450;
  wire net_20452;
  wire net_20453;
  wire net_20455;
  wire net_20459;
  wire net_20460;
  wire net_20466;
  wire net_20470;
  wire net_20471;
  wire net_20472;
  wire net_20476;
  wire net_20477;
  wire net_20478;
  wire net_20483;
  wire net_20484;
  wire net_20489;
  wire net_20490;
  wire net_20495;
  wire net_20496;
  wire net_20501;
  wire net_20502;
  wire net_20507;
  wire net_20508;
  wire net_20513;
  wire net_20514;
  wire net_20517;
  wire net_20519;
  wire net_20520;
  wire net_20527;
  wire net_20531;
  wire net_20532;
  wire net_20533;
  wire net_20535;
  wire net_20536;
  wire net_20538;
  wire net_20552;
  wire net_20560;
  wire net_20566;
  wire net_20584;
  wire net_20591;
  wire net_20593;
  wire net_20596;
  wire net_20598;
  wire net_20601;
  wire net_20602;
  wire net_20606;
  wire net_20611;
  wire net_20625;
  wire net_20629;
  wire net_20637;
  wire net_20644;
  wire net_20647;
  wire net_20652;
  wire net_20653;
  wire net_20655;
  wire net_20656;
  wire net_20657;
  wire net_20658;
  wire net_20659;
  wire net_20660;
  wire net_20661;
  wire net_20695;
  wire net_20712;
  wire net_20713;
  wire net_20715;
  wire net_20717;
  wire net_20721;
  wire net_20725;
  wire net_20726;
  wire net_20728;
  wire net_20737;
  wire net_20743;
  wire net_20746;
  wire net_20752;
  wire net_20759;
  wire net_20766;
  wire net_20770;
  wire net_20775;
  wire net_20776;
  wire net_20779;
  wire net_20782;
  wire net_20783;
  wire net_20784;
  wire net_20806;
  wire net_20818;
  wire net_20825;
  wire net_20831;
  wire net_20834;
  wire net_20841;
  wire net_20846;
  wire net_20852;
  wire net_20858;
  wire net_20877;
  wire net_20883;
  wire net_20888;
  wire net_20896;
  wire net_20898;
  wire net_20899;
  wire net_20901;
  wire net_20930;
  wire net_20942;
  wire net_20949;
  wire net_20952;
  wire net_20954;
  wire net_20955;
  wire net_20958;
  wire net_20967;
  wire net_20977;
  wire net_20980;
  wire net_20993;
  wire net_21001;
  wire net_21006;
  wire net_21013;
  wire net_21017;
  wire net_21021;
  wire net_21022;
  wire net_21024;
  wire net_21026;
  wire net_21027;
  wire net_21035;
  wire net_21038;
  wire net_21045;
  wire net_21070;
  wire net_21075;
  wire net_21078;
  wire net_21088;
  wire net_21091;
  wire net_21115;
  wire net_21116;
  wire net_21117;
  wire net_21118;
  wire net_21143;
  wire net_21144;
  wire net_21145;
  wire net_21146;
  wire net_21150;
  wire net_21161;
  wire net_21192;
  wire net_21196;
  wire net_21205;
  wire net_21222;
  wire net_21258;
  wire net_21264;
  wire net_21267;
  wire net_21268;
  wire net_21280;
  wire net_21315;
  wire net_21317;
  wire net_21368;
  wire net_21375;
  wire net_21390;
  wire net_21391;
  wire net_21579;
  wire net_21626;
  wire net_21636;
  wire net_21637;
  wire net_22622;
  wire net_22697;
  wire net_22721;
  wire net_22746;
  wire net_22756;
  wire net_22785;
  wire net_22790;
  wire net_22791;
  wire net_22815;
  wire net_22817;
  wire net_22818;
  wire net_22841;
  wire net_22844;
  wire net_22845;
  wire net_22846;
  wire net_22848;
  wire net_22861;
  wire net_22874;
  wire net_22895;
  wire net_22898;
  wire net_22944;
  wire net_22955;
  wire net_22968;
  wire net_22990;
  wire net_23006;
  wire net_23007;
  wire net_23013;
  wire net_23014;
  wire net_23015;
  wire net_23016;
  wire net_23055;
  wire net_23056;
  wire net_23061;
  wire net_23063;
  wire net_23069;
  wire net_23071;
  wire net_23077;
  wire net_23078;
  wire net_23095;
  wire net_23108;
  wire net_23113;
  wire net_23125;
  wire net_23126;
  wire net_23127;
  wire net_23128;
  wire net_23129;
  wire net_23130;
  wire net_23132;
  wire net_23133;
  wire net_23134;
  wire net_23135;
  wire net_23136;
  wire net_23137;
  wire net_23138;
  wire net_23139;
  wire net_23157;
  wire net_23177;
  wire net_23179;
  wire net_23186;
  wire net_23188;
  wire net_23189;
  wire net_23190;
  wire net_23197;
  wire net_23198;
  wire net_23204;
  wire net_23206;
  wire net_23215;
  wire net_23220;
  wire net_23224;
  wire net_23225;
  wire net_23232;
  wire net_23237;
  wire net_23243;
  wire net_23251;
  wire net_23253;
  wire net_23254;
  wire net_23266;
  wire net_23273;
  wire net_23283;
  wire net_23286;
  wire net_23287;
  wire net_23288;
  wire net_23289;
  wire net_23299;
  wire net_23301;
  wire net_23305;
  wire net_23306;
  wire net_23307;
  wire net_23308;
  wire net_23310;
  wire net_23327;
  wire net_23328;
  wire net_23330;
  wire net_23331;
  wire net_23334;
  wire net_23336;
  wire net_23338;
  wire net_23340;
  wire net_23342;
  wire net_23344;
  wire net_23346;
  wire net_23348;
  wire net_23350;
  wire net_23352;
  wire net_23354;
  wire net_23356;
  wire net_23358;
  wire net_23361;
  wire net_23362;
  wire net_23364;
  wire net_23366;
  wire net_23368;
  wire net_23374;
  wire net_23376;
  wire net_23377;
  wire net_23389;
  wire net_23390;
  wire net_23391;
  wire net_23392;
  wire net_23402;
  wire net_23419;
  wire net_23421;
  wire net_23422;
  wire net_23423;
  wire net_23424;
  wire net_23425;
  wire net_23426;
  wire net_23427;
  wire net_23436;
  wire net_23443;
  wire net_23445;
  wire net_23446;
  wire net_23448;
  wire net_23451;
  wire net_23453;
  wire net_23454;
  wire net_23457;
  wire net_23459;
  wire net_23460;
  wire net_23461;
  wire net_23463;
  wire net_23465;
  wire net_23466;
  wire net_23467;
  wire net_23469;
  wire net_23471;
  wire net_23472;
  wire net_23473;
  wire net_23475;
  wire net_23477;
  wire net_23478;
  wire net_23479;
  wire net_23481;
  wire net_23483;
  wire net_23484;
  wire net_23485;
  wire net_23491;
  wire net_23496;
  wire net_23498;
  wire net_23499;
  wire net_23515;
  wire net_23517;
  wire net_23536;
  wire net_23547;
  wire net_23548;
  wire net_23551;
  wire net_23553;
  wire net_23554;
  wire net_23555;
  wire net_23556;
  wire net_23567;
  wire net_23571;
  wire net_23581;
  wire net_23582;
  wire net_23583;
  wire net_23584;
  wire net_23589;
  wire net_23593;
  wire net_23594;
  wire net_23595;
  wire net_23605;
  wire net_23606;
  wire net_23607;
  wire net_23608;
  wire net_23621;
  wire net_23622;
  wire net_23636;
  wire net_23640;
  wire net_23668;
  wire net_23670;
  wire net_23671;
  wire net_23672;
  wire net_23674;
  wire net_23676;
  wire net_23678;
  wire net_23682;
  wire net_23684;
  wire net_23687;
  wire net_23700;
  wire net_23704;
  wire net_23706;
  wire net_23711;
  wire net_23716;
  wire net_23719;
  wire net_23722;
  wire net_23728;
  wire net_23736;
  wire net_23741;
  wire net_23745;
  wire net_23746;
  wire net_23747;
  wire net_23748;
  wire net_23749;
  wire net_23750;
  wire net_23751;
  wire net_23752;
  wire net_23753;
  wire net_23754;
  wire net_23767;
  wire net_23769;
  wire net_23771;
  wire net_23773;
  wire net_23774;
  wire net_23775;
  wire net_23778;
  wire net_23779;
  wire net_23781;
  wire net_23782;
  wire net_23804;
  wire net_23805;
  wire net_23806;
  wire net_23807;
  wire net_23811;
  wire net_23812;
  wire net_23814;
  wire net_23817;
  wire net_23822;
  wire net_23828;
  wire net_23834;
  wire net_23842;
  wire net_23848;
  wire net_23851;
  wire net_23860;
  wire net_23866;
  wire net_23868;
  wire net_23869;
  wire net_23870;
  wire net_23871;
  wire net_23872;
  wire net_23873;
  wire net_23874;
  wire net_23875;
  wire net_23876;
  wire net_23877;
  wire net_23882;
  wire net_23905;
  wire net_23914;
  wire net_23916;
  wire net_23918;
  wire net_23920;
  wire net_23929;
  wire net_23933;
  wire net_23937;
  wire net_23939;
  wire net_23947;
  wire net_23953;
  wire net_23956;
  wire net_23964;
  wire net_23968;
  wire net_23974;
  wire net_23981;
  wire net_23986;
  wire net_23990;
  wire net_23991;
  wire net_23993;
  wire net_23994;
  wire net_23995;
  wire net_23996;
  wire net_23997;
  wire net_23998;
  wire net_23999;
  wire net_24000;
  wire net_24006;
  wire net_24007;
  wire net_24020;
  wire net_24024;
  wire net_24042;
  wire net_24049;
  wire net_24050;
  wire net_24052;
  wire net_24054;
  wire net_24058;
  wire net_24060;
  wire net_24062;
  wire net_24067;
  wire net_24074;
  wire net_24081;
  wire net_24087;
  wire net_24092;
  wire net_24098;
  wire net_24104;
  wire net_24109;
  wire net_24114;
  wire net_24115;
  wire net_24116;
  wire net_24117;
  wire net_24118;
  wire net_24119;
  wire net_24120;
  wire net_24121;
  wire net_24122;
  wire net_24123;
  wire net_24136;
  wire net_24145;
  wire net_24146;
  wire net_24147;
  wire net_24148;
  wire net_24161;
  wire net_24164;
  wire net_24170;
  wire net_24173;
  wire net_24175;
  wire net_24177;
  wire net_24182;
  wire net_24184;
  wire net_24193;
  wire net_24199;
  wire net_24202;
  wire net_24211;
  wire net_24216;
  wire net_24221;
  wire net_24226;
  wire net_24235;
  wire net_24237;
  wire net_24238;
  wire net_24256;
  wire net_24263;
  wire net_24265;
  wire net_24268;
  wire net_24283;
  wire net_24286;
  wire net_24293;
  wire net_24296;
  wire net_24298;
  wire net_24300;
  wire net_24306;
  wire net_24310;
  wire net_24313;
  wire net_24320;
  wire net_24328;
  wire net_24333;
  wire net_24337;
  wire net_24344;
  wire net_24350;
  wire net_24358;
  wire net_24360;
  wire net_24361;
  wire net_24392;
  wire net_24416;
  wire net_24421;
  wire net_24423;
  wire net_24428;
  wire net_24431;
  wire net_24432;
  wire net_24438;
  wire net_24443;
  wire net_24451;
  wire net_24462;
  wire net_24469;
  wire net_24479;
  wire net_24483;
  wire net_24484;
  wire net_24512;
  wire net_24533;
  wire net_24535;
  wire net_24538;
  wire net_24548;
  wire net_24551;
  wire net_24553;
  wire net_24557;
  wire net_24566;
  wire net_24571;
  wire net_24578;
  wire net_24583;
  wire net_24590;
  wire net_24598;
  wire net_24601;
  wire net_24606;
  wire net_24607;
  wire net_24634;
  wire net_24639;
  wire net_24649;
  wire net_24651;
  wire net_24653;
  wire net_24654;
  wire net_24656;
  wire net_24657;
  wire net_24658;
  wire net_24659;
  wire net_24660;
  wire net_24661;
  wire net_24662;
  wire net_24665;
  wire net_24675;
  wire net_24676;
  wire net_24680;
  wire net_24694;
  wire net_24695;
  wire net_24696;
  wire net_24697;
  wire net_24712;
  wire net_24713;
  wire net_24714;
  wire net_24715;
  wire net_24718;
  wire net_24719;
  wire net_24720;
  wire net_24721;
  wire net_24724;
  wire net_24725;
  wire net_24726;
  wire net_24727;
  wire net_24728;
  wire net_24729;
  wire net_24730;
  wire net_24772;
  wire net_24773;
  wire net_24780;
  wire net_24783;
  wire net_24792;
  wire net_24811;
  wire net_24812;
  wire net_24813;
  wire net_24814;
  wire net_24851;
  wire net_24852;
  wire net_24853;
  wire net_24870;
  wire net_24895;
  wire net_24899;
  wire net_24925;
  wire net_24937;
  wire net_24948;
  wire net_24952;
  wire net_24974;
  wire net_24975;
  wire net_25024;
  wire net_25038;
  wire net_25053;
  wire net_25077;
  wire net_25098;
  wire net_25099;
  wire net_25111;
  wire net_26358;
  wire net_26453;
  wire net_26489;
  wire net_26554;
  wire net_26631;
  wire net_26632;
  wire net_26633;
  wire net_26721;
  wire net_26767;
  wire net_26769;
  wire net_26770;
  wire net_26771;
  wire net_26839;
  wire net_26841;
  wire net_26843;
  wire net_26844;
  wire net_26847;
  wire net_26849;
  wire net_26850;
  wire net_26853;
  wire net_26855;
  wire net_26856;
  wire net_26860;
  wire net_26861;
  wire net_26862;
  wire net_26866;
  wire net_26867;
  wire net_26869;
  wire net_26870;
  wire net_26871;
  wire net_26872;
  wire net_26874;
  wire net_26876;
  wire net_26877;
  wire net_26878;
  wire net_26879;
  wire net_26880;
  wire net_26881;
  wire net_26882;
  wire net_26883;
  wire net_26884;
  wire net_26885;
  wire net_26886;
  wire net_26888;
  wire net_26889;
  wire net_26890;
  wire net_26891;
  wire net_26896;
  wire net_26897;
  wire net_26898;
  wire net_26899;
  wire net_26900;
  wire net_26905;
  wire net_26906;
  wire net_26914;
  wire net_26939;
  wire net_26943;
  wire net_26944;
  wire net_26945;
  wire net_26949;
  wire net_26950;
  wire net_26951;
  wire net_26952;
  wire net_26955;
  wire net_26956;
  wire net_26957;
  wire net_26960;
  wire net_26961;
  wire net_26962;
  wire net_26964;
  wire net_26965;
  wire net_26968;
  wire net_26969;
  wire net_26972;
  wire net_26973;
  wire net_26974;
  wire net_26975;
  wire net_26976;
  wire net_26977;
  wire net_26978;
  wire net_26979;
  wire net_26980;
  wire net_26981;
  wire net_26982;
  wire net_26983;
  wire net_26984;
  wire net_26985;
  wire net_26986;
  wire net_26987;
  wire net_26988;
  wire net_26990;
  wire net_26991;
  wire net_26992;
  wire net_26993;
  wire net_26998;
  wire net_26999;
  wire net_27000;
  wire net_27001;
  wire net_27002;
  wire net_27003;
  wire net_27004;
  wire net_27005;
  wire net_27006;
  wire net_27007;
  wire net_27008;
  wire net_27025;
  wire net_27028;
  wire net_27032;
  wire net_27074;
  wire net_27075;
  wire net_27076;
  wire net_27077;
  wire net_27078;
  wire net_27079;
  wire net_27080;
  wire net_27118;
  wire net_27135;
  wire net_27175;
  wire net_27176;
  wire net_27177;
  wire net_27178;
  wire net_27179;
  wire net_27180;
  wire net_27181;
  wire net_27182;
  wire net_27235;
  wire net_27277;
  wire net_27278;
  wire net_27279;
  wire net_27280;
  wire net_27281;
  wire net_27282;
  wire net_27283;
  wire net_27284;
  wire net_27338;
  wire net_27379;
  wire net_27380;
  wire net_27381;
  wire net_27382;
  wire net_27383;
  wire net_27385;
  wire net_27386;
  wire net_27435;
  wire net_27444;
  wire net_27467;
  wire net_27469;
  wire net_27471;
  wire net_27477;
  wire net_27481;
  wire net_27482;
  wire net_27483;
  wire net_27484;
  wire net_27485;
  wire net_27487;
  wire net_27488;
  wire net_27497;
  wire net_27498;
  wire net_27508;
  wire net_27509;
  wire net_27510;
  wire net_27524;
  wire net_27535;
  wire net_27537;
  wire net_27569;
  wire net_27583;
  wire net_27584;
  wire net_27585;
  wire net_27586;
  wire net_27587;
  wire net_27588;
  wire net_27589;
  wire net_27590;
  wire net_27610;
  wire net_27611;
  wire net_27627;
  wire net_27635;
  wire net_27640;
  wire net_27647;
  wire net_27655;
  wire net_27657;
  wire net_27659;
  wire net_27665;
  wire net_27686;
  wire net_27687;
  wire net_27688;
  wire net_27689;
  wire net_27690;
  wire net_27691;
  wire net_27692;
  wire net_27701;
  wire net_27702;
  wire net_27712;
  wire net_27713;
  wire net_27714;
  wire net_27731;
  wire net_27738;
  wire net_27739;
  wire net_27743;
  wire net_27746;
  wire net_27766;
  wire net_27787;
  wire net_27788;
  wire net_27789;
  wire net_27790;
  wire net_27791;
  wire net_27792;
  wire net_27793;
  wire net_27794;
  wire net_27814;
  wire net_27815;
  wire net_27844;
  wire net_27850;
  wire net_27892;
  wire net_27893;
  wire net_27895;
  wire net_27896;
  wire net_27943;
  wire net_27947;
  wire net_27991;
  wire net_27992;
  wire net_27993;
  wire net_27994;
  wire net_27995;
  wire net_27996;
  wire net_27997;
  wire net_27998;
  wire net_28036;
  wire net_28093;
  wire net_28095;
  wire net_28096;
  wire net_28097;
  wire net_28100;
  wire net_28136;
  wire net_28202;
  wire net_28297;
  wire net_28299;
  wire net_28300;
  wire net_28301;
  wire net_28302;
  wire net_28303;
  wire net_28399;
  wire net_28402;
  wire net_28404;
  wire net_28405;
  wire net_28542;
  wire net_29689;
  wire net_29728;
  wire net_29752;
  wire net_29755;
  wire net_29756;
  wire net_29758;
  wire net_29759;
  wire net_29760;
  wire net_29823;
  wire net_29834;
  wire net_29875;
  wire net_29876;
  wire net_29881;
  wire net_29883;
  wire net_29887;
  wire net_29961;
  wire net_29980;
  wire net_29983;
  wire net_30003;
  wire net_30010;
  wire net_30018;
  wire net_30038;
  wire net_30039;
  wire net_30040;
  wire net_30045;
  wire net_30046;
  wire net_30047;
  wire net_30069;
  wire net_30081;
  wire net_30091;
  wire net_30104;
  wire net_30112;
  wire net_30116;
  wire net_30126;
  wire net_30132;
  wire net_30139;
  wire net_30161;
  wire net_30162;
  wire net_30163;
  wire net_30165;
  wire net_30166;
  wire net_30167;
  wire net_30168;
  wire net_30169;
  wire net_30170;
  wire net_30175;
  wire net_30182;
  wire net_30185;
  wire net_30189;
  wire net_30208;
  wire net_30211;
  wire net_30221;
  wire net_30224;
  wire net_30225;
  wire net_30232;
  wire net_30235;
  wire net_30237;
  wire net_30244;
  wire net_30252;
  wire net_30255;
  wire net_30268;
  wire net_30269;
  wire net_30281;
  wire net_30284;
  wire net_30285;
  wire net_30286;
  wire net_30287;
  wire net_30288;
  wire net_30289;
  wire net_30290;
  wire net_30291;
  wire net_30292;
  wire net_30293;
  wire net_30296;
  wire net_30301;
  wire net_30302;
  wire net_30305;
  wire net_30308;
  wire net_30310;
  wire net_30320;
  wire net_30321;
  wire net_30329;
  wire net_30333;
  wire net_30336;
  wire net_30337;
  wire net_30341;
  wire net_30342;
  wire net_30343;
  wire net_30346;
  wire net_30348;
  wire net_30350;
  wire net_30354;
  wire net_30355;
  wire net_30358;
  wire net_30359;
  wire net_30361;
  wire net_30362;
  wire net_30365;
  wire net_30367;
  wire net_30368;
  wire net_30369;
  wire net_30371;
  wire net_30373;
  wire net_30374;
  wire net_30375;
  wire net_30378;
  wire net_30380;
  wire net_30381;
  wire net_30385;
  wire net_30386;
  wire net_30387;
  wire net_30392;
  wire net_30393;
  wire net_30396;
  wire net_30397;
  wire net_30398;
  wire net_30399;
  wire net_30403;
  wire net_30406;
  wire net_30407;
  wire net_30409;
  wire net_30410;
  wire net_30412;
  wire net_30413;
  wire net_30414;
  wire net_30415;
  wire net_30416;
  wire net_30420;
  wire net_30423;
  wire net_30436;
  wire net_30440;
  wire net_30442;
  wire net_30453;
  wire net_30455;
  wire net_30459;
  wire net_30460;
  wire net_30461;
  wire net_30463;
  wire net_30476;
  wire net_30477;
  wire net_30478;
  wire net_30481;
  wire net_30482;
  wire net_30484;
  wire net_30485;
  wire net_30488;
  wire net_30490;
  wire net_30491;
  wire net_30492;
  wire net_30494;
  wire net_30496;
  wire net_30497;
  wire net_30498;
  wire net_30501;
  wire net_30502;
  wire net_30504;
  wire net_30508;
  wire net_30516;
  wire net_30521;
  wire net_30525;
  wire net_30526;
  wire net_30530;
  wire net_30531;
  wire net_30532;
  wire net_30534;
  wire net_30538;
  wire net_30560;
  wire net_30564;
  wire net_30565;
  wire net_30575;
  wire net_30576;
  wire net_30579;
  wire net_30580;
  wire net_30584;
  wire net_30591;
  wire net_30592;
  wire net_30601;
  wire net_30604;
  wire net_30608;
  wire net_30614;
  wire net_30621;
  wire net_30625;
  wire net_30630;
  wire net_30632;
  wire net_30636;
  wire net_30639;
  wire net_30645;
  wire net_30649;
  wire net_30653;
  wire net_30654;
  wire net_30656;
  wire net_30657;
  wire net_30658;
  wire net_30659;
  wire net_30660;
  wire net_30661;
  wire net_30662;
  wire net_30696;
  wire net_30702;
  wire net_30704;
  wire net_30712;
  wire net_30718;
  wire net_30720;
  wire net_30724;
  wire net_30726;
  wire net_30732;
  wire net_30735;
  wire net_30743;
  wire net_30747;
  wire net_30755;
  wire net_30760;
  wire net_30766;
  wire net_30774;
  wire net_30776;
  wire net_30777;
  wire net_30778;
  wire net_30779;
  wire net_30780;
  wire net_30782;
  wire net_30783;
  wire net_30784;
  wire net_30785;
  wire net_30793;
  wire net_30798;
  wire net_30813;
  wire net_30820;
  wire net_30828;
  wire net_30830;
  wire net_30831;
  wire net_30836;
  wire net_30841;
  wire net_30848;
  wire net_30852;
  wire net_30861;
  wire net_30865;
  wire net_30873;
  wire net_30876;
  wire net_30891;
  wire net_30896;
  wire net_30898;
  wire net_30899;
  wire net_30902;
  wire net_30903;
  wire net_30927;
  wire net_30936;
  wire net_30946;
  wire net_30950;
  wire net_30958;
  wire net_30959;
  wire net_30963;
  wire net_30967;
  wire net_30969;
  wire net_30975;
  wire net_30983;
  wire net_30988;
  wire net_30993;
  wire net_31001;
  wire net_31011;
  wire net_31018;
  wire net_31022;
  wire net_31023;
  wire net_31024;
  wire net_31025;
  wire net_31026;
  wire net_31027;
  wire net_31028;
  wire net_31029;
  wire net_31030;
  wire net_31031;
  wire net_31048;
  wire net_31051;
  wire net_31053;
  wire net_31054;
  wire net_31071;
  wire net_31076;
  wire net_31079;
  wire net_31084;
  wire net_31086;
  wire net_31087;
  wire net_31091;
  wire net_31095;
  wire net_31100;
  wire net_31104;
  wire net_31111;
  wire net_31117;
  wire net_31123;
  wire net_31128;
  wire net_31134;
  wire net_31140;
  wire net_31145;
  wire net_31146;
  wire net_31154;
  wire net_31164;
  wire net_31165;
  wire net_31169;
  wire net_31172;
  wire net_31177;
  wire net_31179;
  wire net_31189;
  wire net_31190;
  wire net_31191;
  wire net_31192;
  wire net_31195;
  wire net_31196;
  wire net_31197;
  wire net_31198;
  wire net_31199;
  wire net_31201;
  wire net_31203;
  wire net_31207;
  wire net_31214;
  wire net_31217;
  wire net_31220;
  wire net_31222;
  wire net_31223;
  wire net_31226;
  wire net_31228;
  wire net_31229;
  wire net_31230;
  wire net_31232;
  wire net_31234;
  wire net_31235;
  wire net_31236;
  wire net_31238;
  wire net_31240;
  wire net_31241;
  wire net_31242;
  wire net_31244;
  wire net_31246;
  wire net_31247;
  wire net_31248;
  wire net_31250;
  wire net_31252;
  wire net_31253;
  wire net_31254;
  wire net_31256;
  wire net_31258;
  wire net_31259;
  wire net_31260;
  wire net_31266;
  wire net_31270;
  wire net_31271;
  wire net_31272;
  wire net_31273;
  wire net_31274;
  wire net_31275;
  wire net_31276;
  wire net_31277;
  wire net_31300;
  wire net_31304;
  wire net_31312;
  wire net_31313;
  wire net_31314;
  wire net_31315;
  wire net_31319;
  wire net_31322;
  wire net_31331;
  wire net_31340;
  wire net_31344;
  wire net_31353;
  wire net_31356;
  wire net_31364;
  wire net_31368;
  wire net_31376;
  wire net_31382;
  wire net_31386;
  wire net_31391;
  wire net_31392;
  wire net_31393;
  wire net_31399;
  wire net_31444;
  wire net_31445;
  wire net_31448;
  wire net_31459;
  wire net_31486;
  wire net_31494;
  wire net_31505;
  wire net_31511;
  wire net_31514;
  wire net_31515;
  wire net_31516;
  wire net_31517;
  wire net_31518;
  wire net_31519;
  wire net_31520;
  wire net_31522;
  wire net_31523;
  wire net_31532;
  wire net_31546;
  wire net_31557;
  wire net_31558;
  wire net_31559;
  wire net_31561;
  wire net_31562;
  wire net_31563;
  wire net_31564;
  wire net_31565;
  wire net_31566;
  wire net_31567;
  wire net_31568;
  wire net_31569;
  wire net_31570;
  wire net_31571;
  wire net_31572;
  wire net_31573;
  wire net_31574;
  wire net_31575;
  wire net_31577;
  wire net_31578;
  wire net_31582;
  wire net_31583;
  wire net_31584;
  wire net_31585;
  wire net_31586;
  wire net_31590;
  wire net_31591;
  wire net_31592;
  wire net_31593;
  wire net_31596;
  wire net_31597;
  wire net_31598;
  wire net_31599;
  wire net_31602;
  wire net_31603;
  wire net_31604;
  wire net_31605;
  wire net_31608;
  wire net_31609;
  wire net_31610;
  wire net_31611;
  wire net_31614;
  wire net_31615;
  wire net_31616;
  wire net_31617;
  wire net_31620;
  wire net_31621;
  wire net_31622;
  wire net_31623;
  wire net_31628;
  wire net_31632;
  wire net_31633;
  wire net_31634;
  wire net_31635;
  wire net_31636;
  wire net_31637;
  wire net_31638;
  wire net_31640;
  wire net_31642;
  wire net_31645;
  wire net_31652;
  wire net_31696;
  wire net_31699;
  wire net_31701;
  wire net_31709;
  wire net_31711;
  wire net_31716;
  wire net_31727;
  wire net_31731;
  wire net_31737;
  wire net_31756;
  wire net_31760;
  wire net_31761;
  wire net_31805;
  wire net_31806;
  wire net_31807;
  wire net_31808;
  wire net_31811;
  wire net_31812;
  wire net_31813;
  wire net_31814;
  wire net_31816;
  wire net_31817;
  wire net_31818;
  wire net_31824;
  wire net_31832;
  wire net_31833;
  wire net_31837;
  wire net_31838;
  wire net_31843;
  wire net_31844;
  wire net_31849;
  wire net_31850;
  wire net_31855;
  wire net_31856;
  wire net_31861;
  wire net_31862;
  wire net_31867;
  wire net_31868;
  wire net_31871;
  wire net_31873;
  wire net_31874;
  wire net_31881;
  wire net_31883;
  wire net_31884;
  wire net_31932;
  wire net_31934;
  wire net_31937;
  wire net_31939;
  wire net_31954;
  wire net_31956;
  wire net_31961;
  wire net_31971;
  wire net_31979;
  wire net_31986;
  wire net_31991;
  wire net_31995;
  wire net_32006;
  wire net_32007;
  wire net_32065;
  wire net_32070;
  wire net_32072;
  wire net_32074;
  wire net_32084;
  wire net_32102;
  wire net_32113;
  wire net_32119;
  wire net_32129;
  wire net_32130;
  wire net_33484;
  wire net_33486;
  wire net_33559;
  wire net_33572;
  wire net_33585;
  wire net_33587;
  wire net_33588;
  wire net_33590;
  wire net_33591;
  wire net_33605;
  wire net_33635;
  wire net_33644;
  wire net_33646;
  wire net_33648;
  wire net_33652;
  wire net_33673;
  wire net_33678;
  wire net_33689;
  wire net_33695;
  wire net_33704;
  wire net_33706;
  wire net_33707;
  wire net_33715;
  wire net_33718;
  wire net_33771;
  wire net_33812;
  wire net_33813;
  wire net_33818;
  wire net_33824;
  wire net_33835;
  wire net_33859;
  wire net_33869;
  wire net_33870;
  wire net_33874;
  wire net_33877;
  wire net_33889;
  wire net_33896;
  wire net_33900;
  wire net_33904;
  wire net_33914;
  wire net_33917;
  wire net_33918;
  wire net_33931;
  wire net_33933;
  wire net_33934;
  wire net_33935;
  wire net_33937;
  wire net_33941;
  wire net_33945;
  wire net_33946;
  wire net_33947;
  wire net_33948;
  wire net_33975;
  wire net_33981;
  wire net_33982;
  wire net_33983;
  wire net_33984;
  wire net_33990;
  wire net_33991;
  wire net_33992;
  wire net_33994;
  wire net_33996;
  wire net_33999;
  wire net_34000;
  wire net_34001;
  wire net_34038;
  wire net_34040;
  wire net_34045;
  wire net_34053;
  wire net_34055;
  wire net_34056;
  wire net_34064;
  wire net_34071;
  wire net_34080;
  wire net_34086;
  wire net_34092;
  wire net_34099;
  wire net_34107;
  wire net_34110;
  wire net_34115;
  wire net_34116;
  wire net_34117;
  wire net_34118;
  wire net_34120;
  wire net_34121;
  wire net_34123;
  wire net_34124;
  wire net_34126;
  wire net_34148;
  wire net_34152;
  wire net_34160;
  wire net_34167;
  wire net_34171;
  wire net_34179;
  wire net_34181;
  wire net_34185;
  wire net_34186;
  wire net_34187;
  wire net_34189;
  wire net_34192;
  wire net_34197;
  wire net_34205;
  wire net_34212;
  wire net_34215;
  wire net_34217;
  wire net_34222;
  wire net_34224;
  wire net_34227;
  wire net_34235;
  wire net_34238;
  wire net_34239;
  wire net_34240;
  wire net_34242;
  wire net_34243;
  wire net_34244;
  wire net_34251;
  wire net_34252;
  wire net_34284;
  wire net_34286;
  wire net_34294;
  wire net_34298;
  wire net_34300;
  wire net_34304;
  wire net_34306;
  wire net_34314;
  wire net_34323;
  wire net_34332;
  wire net_34341;
  wire net_34346;
  wire net_34353;
  wire net_34356;
  wire net_34360;
  wire net_34361;
  wire net_34363;
  wire net_34364;
  wire net_34365;
  wire net_34366;
  wire net_34367;
  wire net_34368;
  wire net_34369;
  wire net_34370;
  wire net_34375;
  wire net_34378;
  wire net_34387;
  wire net_34389;
  wire net_34391;
  wire net_34406;
  wire net_34409;
  wire net_34418;
  wire net_34439;
  wire net_34450;
  wire net_34476;
  wire net_34483;
  wire net_34484;
  wire net_34487;
  wire net_34488;
  wire net_34489;
  wire net_34490;
  wire net_34491;
  wire net_34492;
  wire net_34493;
  wire net_34498;
  wire net_34507;
  wire net_34510;
  wire net_34511;
  wire net_34528;
  wire net_34529;
  wire net_34531;
  wire net_34532;
  wire net_34534;
  wire net_34539;
  wire net_34540;
  wire net_34541;
  wire net_34542;
  wire net_34544;
  wire net_34547;
  wire net_34552;
  wire net_34553;
  wire net_34558;
  wire net_34559;
  wire net_34561;
  wire net_34562;
  wire net_34565;
  wire net_34567;
  wire net_34568;
  wire net_34569;
  wire net_34571;
  wire net_34573;
  wire net_34574;
  wire net_34575;
  wire net_34577;
  wire net_34579;
  wire net_34580;
  wire net_34581;
  wire net_34583;
  wire net_34585;
  wire net_34586;
  wire net_34587;
  wire net_34589;
  wire net_34591;
  wire net_34592;
  wire net_34593;
  wire net_34595;
  wire net_34597;
  wire net_34598;
  wire net_34599;
  wire net_34605;
  wire net_34609;
  wire net_34610;
  wire net_34611;
  wire net_34612;
  wire net_34613;
  wire net_34614;
  wire net_34615;
  wire net_34616;
  wire net_34624;
  wire net_34626;
  wire net_34630;
  wire net_34632;
  wire net_34634;
  wire net_34640;
  wire net_34652;
  wire net_34662;
  wire net_34664;
  wire net_34665;
  wire net_34668;
  wire net_34672;
  wire net_34676;
  wire net_34678;
  wire net_34686;
  wire net_34691;
  wire net_34692;
  wire net_34696;
  wire net_34709;
  wire net_34714;
  wire net_34722;
  wire net_34726;
  wire net_34730;
  wire net_34731;
  wire net_34732;
  wire net_34733;
  wire net_34734;
  wire net_34736;
  wire net_34737;
  wire net_34738;
  wire net_34739;
  wire net_34756;
  wire net_34759;
  wire net_34760;
  wire net_34773;
  wire net_34788;
  wire net_34791;
  wire net_34813;
  wire net_34820;
  wire net_34852;
  wire net_34853;
  wire net_34855;
  wire net_34861;
  wire net_34873;
  wire net_34877;
  wire net_34882;
  wire net_34884;
  wire net_34889;
  wire net_34904;
  wire net_34906;
  wire net_34908;
  wire net_34916;
  wire net_34918;
  wire net_34920;
  wire net_34922;
  wire net_34926;
  wire net_34932;
  wire net_34937;
  wire net_34942;
  wire net_34947;
  wire net_34953;
  wire net_34962;
  wire net_34968;
  wire net_34971;
  wire net_34976;
  wire net_34977;
  wire net_34978;
  wire net_34979;
  wire net_34982;
  wire net_34983;
  wire net_34990;
  wire net_34991;
  wire net_34997;
  wire net_34998;
  wire net_35010;
  wire net_35021;
  wire net_35023;
  wire net_35028;
  wire net_35030;
  wire net_35032;
  wire net_35033;
  wire net_35034;
  wire net_35035;
  wire net_35040;
  wire net_35053;
  wire net_35054;
  wire net_35059;
  wire net_35066;
  wire net_35071;
  wire net_35078;
  wire net_35083;
  wire net_35087;
  wire net_35089;
  wire net_35093;
  wire net_35095;
  wire net_35097;
  wire net_35099;
  wire net_35100;
  wire net_35104;
  wire net_35106;
  wire net_35107;
  wire net_35120;
  wire net_35122;
  wire net_35127;
  wire net_35129;
  wire net_35130;
  wire net_35131;
  wire net_35137;
  wire net_35154;
  wire net_35158;
  wire net_35161;
  wire net_35168;
  wire net_35170;
  wire net_35172;
  wire net_35173;
  wire net_35178;
  wire net_35181;
  wire net_35189;
  wire net_35193;
  wire net_35202;
  wire net_35207;
  wire net_35212;
  wire net_35218;
  wire net_35222;
  wire net_35223;
  wire net_35224;
  wire net_35226;
  wire net_35227;
  wire net_35228;
  wire net_35229;
  wire net_35231;
  wire net_35232;
  wire net_35251;
  wire net_35254;
  wire net_35269;
  wire net_35273;
  wire net_35276;
  wire net_35281;
  wire net_35282;
  wire net_35298;
  wire net_35334;
  wire net_35335;
  wire net_35336;
  wire net_35337;
  wire net_35344;
  wire net_35345;
  wire net_35347;
  wire net_35348;
  wire net_35349;
  wire net_35350;
  wire net_35351;
  wire net_35352;
  wire net_35353;
  wire net_35354;
  wire net_35359;
  wire net_35368;
  wire net_35372;
  wire net_35378;
  wire net_35388;
  wire net_35390;
  wire net_35391;
  wire net_35392;
  wire net_35394;
  wire net_35396;
  wire net_35397;
  wire net_35399;
  wire net_35400;
  wire net_35401;
  wire net_35402;
  wire net_35403;
  wire net_35404;
  wire net_35405;
  wire net_35406;
  wire net_35407;
  wire net_35410;
  wire net_35413;
  wire net_35414;
  wire net_35415;
  wire net_35416;
  wire net_35417;
  wire net_35419;
  wire net_35421;
  wire net_35422;
  wire net_35423;
  wire net_35424;
  wire net_35427;
  wire net_35428;
  wire net_35429;
  wire net_35430;
  wire net_35433;
  wire net_35434;
  wire net_35435;
  wire net_35436;
  wire net_35439;
  wire net_35440;
  wire net_35441;
  wire net_35442;
  wire net_35445;
  wire net_35446;
  wire net_35447;
  wire net_35448;
  wire net_35457;
  wire net_35458;
  wire net_35459;
  wire net_35460;
  wire net_35463;
  wire net_35464;
  wire net_35465;
  wire net_35466;
  wire net_35467;
  wire net_35468;
  wire net_35470;
  wire net_35473;
  wire net_35474;
  wire net_35475;
  wire net_35477;
  wire net_35482;
  wire net_35485;
  wire net_35488;
  wire net_35497;
  wire net_35499;
  wire net_35513;
  wire net_35515;
  wire net_35519;
  wire net_35522;
  wire net_35524;
  wire net_35525;
  wire net_35526;
  wire net_35528;
  wire net_35530;
  wire net_35533;
  wire net_35535;
  wire net_35536;
  wire net_35550;
  wire net_35551;
  wire net_35552;
  wire net_35553;
  wire net_35562;
  wire net_35563;
  wire net_35564;
  wire net_35565;
  wire net_35580;
  wire net_35581;
  wire net_35582;
  wire net_35583;
  wire net_35590;
  wire net_35591;
  wire net_35592;
  wire net_35593;
  wire net_35594;
  wire net_35595;
  wire net_35596;
  wire net_35619;
  wire net_35716;
  wire net_35717;
  wire net_35718;
  wire net_35721;
  wire net_35722;
  wire net_35723;
  wire net_35973;
  wire net_36219;
  wire net_37390;
  wire net_37393;
  wire net_37403;
  wire net_37406;
  wire net_37416;
  wire net_37417;
  wire net_37420;
  wire net_37421;
  wire net_37422;
  wire net_37438;
  wire net_37457;
  wire net_37462;
  wire net_37464;
  wire net_37468;
  wire net_37480;
  wire net_37498;
  wire net_37510;
  wire net_37516;
  wire net_37529;
  wire net_37533;
  wire net_37537;
  wire net_37538;
  wire net_37543;
  wire net_37544;
  wire net_37545;
  wire net_37546;
  wire net_37547;
  wire net_37548;
  wire net_37549;
  wire net_37550;
  wire net_37597;
  wire net_37631;
  wire net_37633;
  wire net_37672;
  wire net_37691;
  wire net_37699;
  wire net_37700;
  wire net_37702;
  wire net_37703;
  wire net_37704;
  wire net_37705;
  wire net_37706;
  wire net_37707;
  wire net_37708;
  wire net_37709;
  wire net_37716;
  wire net_37719;
  wire net_37720;
  wire net_37729;
  wire net_37743;
  wire net_37746;
  wire net_37749;
  wire net_37752;
  wire net_37754;
  wire net_37762;
  wire net_37795;
  wire net_37812;
  wire net_37813;
  wire net_37814;
  wire net_37815;
  wire net_37822;
  wire net_37823;
  wire net_37825;
  wire net_37826;
  wire net_37828;
  wire net_37830;
  wire net_37831;
  wire net_37832;
  wire net_37844;
  wire net_37849;
  wire net_37857;
  wire net_37868;
  wire net_37870;
  wire net_37872;
  wire net_37873;
  wire net_37876;
  wire net_37880;
  wire net_37884;
  wire net_37885;
  wire net_37895;
  wire net_37899;
  wire net_37900;
  wire net_37901;
  wire net_37902;
  wire net_37914;
  wire net_37929;
  wire net_37937;
  wire net_37942;
  wire net_37945;
  wire net_37946;
  wire net_37949;
  wire net_37952;
  wire net_37953;
  wire net_37954;
  wire net_37955;
  wire net_37966;
  wire net_37974;
  wire net_37983;
  wire net_37989;
  wire net_37995;
  wire net_37997;
  wire net_37998;
  wire net_38008;
  wire net_38011;
  wire net_38016;
  wire net_38024;
  wire net_38031;
  wire net_38040;
  wire net_38041;
  wire net_38047;
  wire net_38058;
  wire net_38060;
  wire net_38065;
  wire net_38069;
  wire net_38070;
  wire net_38072;
  wire net_38075;
  wire net_38078;
  wire net_38087;
  wire net_38102;
  wire net_38118;
  wire net_38119;
  wire net_38120;
  wire net_38127;
  wire net_38145;
  wire net_38160;
  wire net_38166;
  wire net_38172;
  wire net_38192;
  wire net_38193;
  wire net_38194;
  wire net_38195;
  wire net_38197;
  wire net_38198;
  wire net_38199;
  wire net_38201;
  wire net_38213;
  wire net_38219;
  wire net_38228;
  wire net_38236;
  wire net_38240;
  wire net_38242;
  wire net_38244;
  wire net_38246;
  wire net_38249;
  wire net_38253;
  wire net_38255;
  wire net_38256;
  wire net_38269;
  wire net_38276;
  wire net_38280;
  wire net_38286;
  wire net_38294;
  wire net_38298;
  wire net_38299;
  wire net_38304;
  wire net_38312;
  wire net_38315;
  wire net_38316;
  wire net_38317;
  wire net_38318;
  wire net_38320;
  wire net_38321;
  wire net_38322;
  wire net_38323;
  wire net_38324;
  wire net_38326;
  wire net_38336;
  wire net_38346;
  wire net_38359;
  wire net_38361;
  wire net_38363;
  wire net_38364;
  wire net_38365;
  wire net_38368;
  wire net_38370;
  wire net_38373;
  wire net_38375;
  wire net_38380;
  wire net_38390;
  wire net_38392;
  wire net_38393;
  wire net_38396;
  wire net_38398;
  wire net_38399;
  wire net_38400;
  wire net_38402;
  wire net_38404;
  wire net_38406;
  wire net_38408;
  wire net_38411;
  wire net_38412;
  wire net_38414;
  wire net_38416;
  wire net_38418;
  wire net_38420;
  wire net_38423;
  wire net_38424;
  wire net_38426;
  wire net_38429;
  wire net_38430;
  wire net_38432;
  wire net_38435;
  wire net_38436;
  wire net_38438;
  wire net_38439;
  wire net_38443;
  wire net_38457;
  wire net_38464;
  wire net_38466;
  wire net_38476;
  wire net_38484;
  wire net_38485;
  wire net_38486;
  wire net_38487;
  wire net_38491;
  wire net_38494;
  wire net_38495;
  wire net_38517;
  wire net_38522;
  wire net_38528;
  wire net_38532;
  wire net_38539;
  wire net_38544;
  wire net_38550;
  wire net_38559;
  wire net_38561;
  wire net_38562;
  wire net_38563;
  wire net_38564;
  wire net_38565;
  wire net_38566;
  wire net_38568;
  wire net_38569;
  wire net_38570;
  wire net_38588;
  wire net_38592;
  wire net_38593;
  wire net_38596;
  wire net_38604;
  wire net_38608;
  wire net_38614;
  wire net_38615;
  wire net_38616;
  wire net_38624;
  wire net_38629;
  wire net_38632;
  wire net_38639;
  wire net_38643;
  wire net_38649;
  wire net_38662;
  wire net_38670;
  wire net_38675;
  wire net_38679;
  wire net_38680;
  wire net_38684;
  wire net_38685;
  wire net_38686;
  wire net_38687;
  wire net_38689;
  wire net_38690;
  wire net_38692;
  wire net_38693;
  wire net_38701;
  wire net_38703;
  wire net_38720;
  wire net_38735;
  wire net_38738;
  wire net_38749;
  wire net_38760;
  wire net_38761;
  wire net_38796;
  wire net_38797;
  wire net_38806;
  wire net_38807;
  wire net_38808;
  wire net_38811;
  wire net_38852;
  wire net_38858;
  wire net_38873;
  wire net_38877;
  wire net_38879;
  wire net_38880;
  wire net_38886;
  wire net_38891;
  wire net_38908;
  wire net_38914;
  wire net_38916;
  wire net_38929;
  wire net_38930;
  wire net_38933;
  wire net_38934;
  wire net_38955;
  wire net_38958;
  wire net_38982;
  wire net_38983;
  wire net_38984;
  wire net_38990;
  wire net_38991;
  wire net_39000;
  wire net_39003;
  wire net_39026;
  wire net_39039;
  wire net_39042;
  wire net_39043;
  wire net_39044;
  wire net_39045;
  wire net_39052;
  wire net_39053;
  wire net_39055;
  wire net_39056;
  wire net_39058;
  wire net_39059;
  wire net_39060;
  wire net_39062;
  wire net_39068;
  wire net_39069;
  wire net_39098;
  wire net_39099;
  wire net_39100;
  wire net_39107;
  wire net_39110;
  wire net_39114;
  wire net_39115;
  wire net_39118;
  wire net_39123;
  wire net_39126;
  wire net_39129;
  wire net_39130;
  wire net_39131;
  wire net_39132;
  wire net_39141;
  wire net_39148;
  wire net_39156;
  wire net_39162;
  wire net_39171;
  wire net_39175;
  wire net_39176;
  wire net_39178;
  wire net_39180;
  wire net_39182;
  wire net_39185;
  wire net_39197;
  wire net_39224;
  wire net_39228;
  wire net_39230;
  wire net_39231;
  wire net_39233;
  wire net_39234;
  wire net_39235;
  wire net_39236;
  wire net_39238;
  wire net_39244;
  wire net_39246;
  wire net_39247;
  wire net_39249;
  wire net_39254;
  wire net_39258;
  wire net_39259;
  wire net_39260;
  wire net_39261;
  wire net_39266;
  wire net_39272;
  wire net_39276;
  wire net_39277;
  wire net_39278;
  wire net_39279;
  wire net_39284;
  wire net_39291;
  wire net_39294;
  wire net_39298;
  wire net_39299;
  wire net_39301;
  wire net_39302;
  wire net_39304;
  wire net_39305;
  wire net_39306;
  wire net_39314;
  wire net_39318;
  wire net_39325;
  wire net_39331;
  wire net_39344;
  wire net_39345;
  wire net_39348;
  wire net_39352;
  wire net_39360;
  wire net_39364;
  wire net_39376;
  wire net_39394;
  wire net_39401;
  wire net_39406;
  wire net_39419;
  wire net_39421;
  wire net_39422;
  wire net_39424;
  wire net_39425;
  wire net_39426;
  wire net_39428;
  wire net_39430;
  wire net_39431;
  wire net_39436;
  wire net_39453;
  wire net_39455;
  wire net_39458;
  wire net_39466;
  wire net_39474;
  wire net_39476;
  wire net_39480;
  wire net_39481;
  wire net_39482;
  wire net_39483;
  wire net_39484;
  wire net_39492;
  wire net_39498;
  wire net_39504;
  wire net_39505;
  wire net_39506;
  wire net_39507;
  wire net_39510;
  wire net_39511;
  wire net_39512;
  wire net_39513;
  wire net_39518;
  wire net_39544;
  wire net_39545;
  wire net_39547;
  wire net_39548;
  wire net_39549;
  wire net_39550;
  wire net_39551;
  wire net_39552;
  wire net_39553;
  wire net_39554;
  wire net_39581;
  wire net_39588;
  wire net_39589;
  wire net_39590;
  wire net_39591;
  wire net_39592;
  wire net_39594;
  wire net_39595;
  wire net_39596;
  wire net_39597;
  wire net_39598;
  wire net_39599;
  wire net_39600;
  wire net_39602;
  wire net_39603;
  wire net_39604;
  wire net_39608;
  wire net_39610;
  wire net_39612;
  wire net_39613;
  wire net_39615;
  wire net_39618;
  wire net_39621;
  wire net_39622;
  wire net_39623;
  wire net_39624;
  wire net_39627;
  wire net_39628;
  wire net_39629;
  wire net_39630;
  wire net_39633;
  wire net_39634;
  wire net_39635;
  wire net_39636;
  wire net_39651;
  wire net_39652;
  wire net_39653;
  wire net_39654;
  wire net_39657;
  wire net_39658;
  wire net_39659;
  wire net_39660;
  wire net_39663;
  wire net_39664;
  wire net_39665;
  wire net_39666;
  wire net_39667;
  wire net_39668;
  wire net_39671;
  wire net_39677;
  wire net_41250;
  wire net_41270;
  wire net_41289;
  wire net_41292;
  wire net_41293;
  wire net_41294;
  wire net_41299;
  wire net_41302;
  wire net_41303;
  wire net_41309;
  wire net_41320;
  wire net_41322;
  wire net_41323;
  wire net_41326;
  wire net_41328;
  wire net_41329;
  wire net_41330;
  wire net_41333;
  wire net_41334;
  wire net_41336;
  wire net_41352;
  wire net_41358;
  wire net_41365;
  wire net_41366;
  wire net_41368;
  wire net_41369;
  wire net_41375;
  wire net_41376;
  wire net_41378;
  wire net_41379;
  wire net_41380;
  wire net_41381;
  wire net_41397;
  wire net_41431;
  wire net_41440;
  wire net_41452;
  wire net_41457;
  wire net_41458;
  wire net_41470;
  wire net_41474;
  wire net_41475;
  wire net_41477;
  wire net_41479;
  wire net_41485;
  wire net_41490;
  wire net_41497;
  wire net_41504;
  wire net_41511;
  wire net_41517;
  wire net_41521;
  wire net_41526;
  wire net_41531;
  wire net_41532;
  wire net_41534;
  wire net_41535;
  wire net_41536;
  wire net_41537;
  wire net_41538;
  wire net_41539;
  wire net_41540;
  wire net_41558;
  wire net_41559;
  wire net_41560;
  wire net_41564;
  wire net_41566;
  wire net_41584;
  wire net_41589;
  wire net_41593;
  wire net_41594;
  wire net_41595;
  wire net_41598;
  wire net_41603;
  wire net_41604;
  wire net_41608;
  wire net_41615;
  wire net_41622;
  wire net_41627;
  wire net_41633;
  wire net_41637;
  wire net_41645;
  wire net_41650;
  wire net_41654;
  wire net_41655;
  wire net_41657;
  wire net_41658;
  wire net_41659;
  wire net_41660;
  wire net_41661;
  wire net_41662;
  wire net_41663;
  wire net_41668;
  wire net_41674;
  wire net_41682;
  wire net_41686;
  wire net_41688;
  wire net_41703;
  wire net_41704;
  wire net_41706;
  wire net_41708;
  wire net_41710;
  wire net_41712;
  wire net_41714;
  wire net_41719;
  wire net_41724;
  wire net_41725;
  wire net_41727;
  wire net_41730;
  wire net_41731;
  wire net_41732;
  wire net_41733;
  wire net_41737;
  wire net_41750;
  wire net_41761;
  wire net_41766;
  wire net_41772;
  wire net_41773;
  wire net_41774;
  wire net_41775;
  wire net_41776;
  wire net_41777;
  wire net_41779;
  wire net_41780;
  wire net_41781;
  wire net_41782;
  wire net_41783;
  wire net_41784;
  wire net_41785;
  wire net_41786;
  wire net_41792;
  wire net_41793;
  wire net_41796;
  wire net_41828;
  wire net_41832;
  wire net_41842;
  wire net_41846;
  wire net_41849;
  wire net_41859;
  wire net_41877;
  wire net_41886;
  wire net_41892;
  wire net_41895;
  wire net_41900;
  wire net_41901;
  wire net_41902;
  wire net_41903;
  wire net_41906;
  wire net_41909;
  wire net_41926;
  wire net_41931;
  wire net_41953;
  wire net_41960;
  wire net_41968;
  wire net_41983;
  wire net_42001;
  wire net_42018;
  wire net_42022;
  wire net_42023;
  wire net_42025;
  wire net_42029;
  wire net_42030;
  wire net_42041;
  wire net_42046;
  wire net_42048;
  wire net_42057;
  wire net_42070;
  wire net_42072;
  wire net_42073;
  wire net_42074;
  wire net_42082;
  wire net_42091;
  wire net_42093;
  wire net_42100;
  wire net_42107;
  wire net_42118;
  wire net_42123;
  wire net_42125;
  wire net_42130;
  wire net_42144;
  wire net_42146;
  wire net_42147;
  wire net_42148;
  wire net_42149;
  wire net_42150;
  wire net_42151;
  wire net_42152;
  wire net_42153;
  wire net_42154;
  wire net_42155;
  wire net_42156;
  wire net_42160;
  wire net_42193;
  wire net_42198;
  wire net_42199;
  wire net_42202;
  wire net_42203;
  wire net_42213;
  wire net_42218;
  wire net_42225;
  wire net_42229;
  wire net_42240;
  wire net_42248;
  wire net_42255;
  wire net_42259;
  wire net_42265;
  wire net_42269;
  wire net_42270;
  wire net_42272;
  wire net_42275;
  wire net_42278;
  wire net_42281;
  wire net_42294;
  wire net_42296;
  wire net_42302;
  wire net_42306;
  wire net_42319;
  wire net_42365;
  wire net_42391;
  wire net_42392;
  wire net_42395;
  wire net_42398;
  wire net_42401;
  wire net_42402;
  wire net_42412;
  wire net_42416;
  wire net_42436;
  wire net_42437;
  wire net_42439;
  wire net_42444;
  wire net_42445;
  wire net_42448;
  wire net_42454;
  wire net_42456;
  wire net_42470;
  wire net_42475;
  wire net_42480;
  wire net_42486;
  wire net_42500;
  wire net_42505;
  wire net_42506;
  wire net_42512;
  wire net_42515;
  wire net_42516;
  wire net_42517;
  wire net_42518;
  wire net_42519;
  wire net_42520;
  wire net_42521;
  wire net_42522;
  wire net_42523;
  wire net_42524;
  wire net_42526;
  wire net_42529;
  wire net_42558;
  wire net_42559;
  wire net_42560;
  wire net_42565;
  wire net_42567;
  wire net_42569;
  wire net_42572;
  wire net_42575;
  wire net_42576;
  wire net_42581;
  wire net_42588;
  wire net_42594;
  wire net_42598;
  wire net_42609;
  wire net_42615;
  wire net_42616;
  wire net_42617;
  wire net_42618;
  wire net_42630;
  wire net_42633;
  wire net_42634;
  wire net_42635;
  wire net_42636;
  wire net_42637;
  wire net_42638;
  wire net_42640;
  wire net_42641;
  wire net_42642;
  wire net_42644;
  wire net_42645;
  wire net_42659;
  wire net_42672;
  wire net_42683;
  wire net_42692;
  wire net_42726;
  wire net_42760;
  wire net_42761;
  wire net_42765;
  wire net_42767;
  wire net_42791;
  wire net_42794;
  wire net_42798;
  wire net_42806;
  wire net_42810;
  wire net_42814;
  wire net_42843;
  wire net_42851;
  wire net_42883;
  wire net_42884;
  wire net_42886;
  wire net_42888;
  wire net_42890;
  wire net_42891;
  wire net_42893;
  wire net_42927;
  wire net_42936;
  wire net_42951;
  wire net_42952;
  wire net_42953;
  wire net_42954;
  wire net_42955;
  wire net_42961;
  wire net_42969;
  wire net_42980;
  wire net_42985;
  wire net_42993;
  wire net_43003;
  wire net_43006;
  wire net_43007;
  wire net_43009;
  wire net_43010;
  wire net_43011;
  wire net_43013;
  wire net_43015;
  wire net_43016;
  wire net_43023;
  wire net_43028;
  wire net_43034;
  wire net_43044;
  wire net_43052;
  wire net_43053;
  wire net_43056;
  wire net_43061;
  wire net_43063;
  wire net_43065;
  wire net_43076;
  wire net_43077;
  wire net_43085;
  wire net_43095;
  wire net_43096;
  wire net_43097;
  wire net_43098;
  wire net_43109;
  wire net_43128;
  wire net_43129;
  wire net_43130;
  wire net_43132;
  wire net_43133;
  wire net_43135;
  wire net_43136;
  wire net_43146;
  wire net_43152;
  wire net_43156;
  wire net_43165;
  wire net_43182;
  wire net_43187;
  wire net_43191;
  wire net_43192;
  wire net_43193;
  wire net_43196;
  wire net_43207;
  wire net_43215;
  wire net_43226;
  wire net_43231;
  wire net_43237;
  wire net_43252;
  wire net_43253;
  wire net_43255;
  wire net_43257;
  wire net_43258;
  wire net_43259;
  wire net_43260;
  wire net_43261;
  wire net_43262;
  wire net_43272;
  wire net_43276;
  wire net_43281;
  wire net_43296;
  wire net_43298;
  wire net_43299;
  wire net_43300;
  wire net_43301;
  wire net_43302;
  wire net_43305;
  wire net_43307;
  wire net_43310;
  wire net_43315;
  wire net_43316;
  wire net_43319;
  wire net_43329;
  wire net_43330;
  wire net_43331;
  wire net_43332;
  wire net_43335;
  wire net_43341;
  wire net_43342;
  wire net_43343;
  wire net_43344;
  wire net_43353;
  wire net_43365;
  wire net_43366;
  wire net_43367;
  wire net_43368;
  wire net_43372;
  wire net_43375;
  wire net_43376;
  wire net_43379;
  wire net_43380;
  wire net_43383;
  wire net_43385;
  wire net_43393;
  wire net_43405;
  wire net_43419;
  wire net_43421;
  wire net_43422;
  wire net_43425;
  wire net_43426;
  wire net_43428;
  wire net_43431;
  wire net_43432;
  wire net_43434;
  wire net_43435;
  wire net_43437;
  wire net_43438;
  wire net_43439;
  wire net_43441;
  wire net_43444;
  wire net_43448;
  wire net_43450;
  wire net_43452;
  wire net_43453;
  wire net_43454;
  wire net_43458;
  wire net_43459;
  wire net_43460;
  wire net_43465;
  wire net_43466;
  wire net_43467;
  wire net_43470;
  wire net_43471;
  wire net_43473;
  wire net_43476;
  wire net_43477;
  wire net_43478;
  wire net_43483;
  wire net_43484;
  wire net_43485;
  wire net_43488;
  wire net_43489;
  wire net_43491;
  wire net_43495;
  wire net_43496;
  wire net_43497;
  wire net_43498;
  wire net_43499;
  wire net_43500;
  wire net_43502;
  wire net_43513;
  wire net_43518;
  wire net_43523;
  wire net_43544;
  wire net_43549;
  wire net_43551;
  wire net_43556;
  wire net_43557;
  wire net_43559;
  wire net_43568;
  wire net_43569;
  wire net_43581;
  wire net_43582;
  wire net_43583;
  wire net_43584;
  wire net_43617;
  wire net_43618;
  wire net_43619;
  wire net_43620;
  wire net_43621;
  wire net_43622;
  wire net_43623;
  wire net_45078;
  wire net_45079;
  wire net_45080;
  wire net_45081;
  wire net_45135;
  wire net_45178;
  wire net_45199;
  wire net_45200;
  wire net_45205;
  wire net_45206;
  wire net_45207;
  wire net_45208;
  wire net_45209;
  wire net_45211;
  wire net_45215;
  wire net_45216;
  wire net_45228;
  wire net_45257;
  wire net_45258;
  wire net_45259;
  wire net_45264;
  wire net_45271;
  wire net_45276;
  wire net_45283;
  wire net_45296;
  wire net_45299;
  wire net_45300;
  wire net_45301;
  wire net_45304;
  wire net_45305;
  wire net_45308;
  wire net_45311;
  wire net_45312;
  wire net_45313;
  wire net_45314;
  wire net_45316;
  wire net_45317;
  wire net_45320;
  wire net_45322;
  wire net_45323;
  wire net_45324;
  wire net_45328;
  wire net_45329;
  wire net_45330;
  wire net_45340;
  wire net_45345;
  wire net_45347;
  wire net_45353;
  wire net_45357;
  wire net_45362;
  wire net_45363;
  wire net_45368;
  wire net_45369;
  wire net_45370;
  wire net_45371;
  wire net_45378;
  wire net_45389;
  wire net_45390;
  wire net_45392;
  wire net_45395;
  wire net_45408;
  wire net_45411;
  wire net_45412;
  wire net_45413;
  wire net_45414;
  wire net_45415;
  wire net_45417;
  wire net_45418;
  wire net_45420;
  wire net_45425;
  wire net_45427;
  wire net_45429;
  wire net_45430;
  wire net_45435;
  wire net_45437;
  wire net_45439;
  wire net_45440;
  wire net_45443;
  wire net_45445;
  wire net_45446;
  wire net_45447;
  wire net_45449;
  wire net_45451;
  wire net_45452;
  wire net_45453;
  wire net_45455;
  wire net_45457;
  wire net_45458;
  wire net_45459;
  wire net_45461;
  wire net_45463;
  wire net_45464;
  wire net_45465;
  wire net_45467;
  wire net_45469;
  wire net_45470;
  wire net_45471;
  wire net_45473;
  wire net_45475;
  wire net_45476;
  wire net_45477;
  wire net_45483;
  wire net_45487;
  wire net_45488;
  wire net_45489;
  wire net_45490;
  wire net_45491;
  wire net_45492;
  wire net_45493;
  wire net_45494;
  wire net_45515;
  wire net_45529;
  wire net_45532;
  wire net_45533;
  wire net_45534;
  wire net_45538;
  wire net_45539;
  wire net_45541;
  wire net_45542;
  wire net_45543;
  wire net_45546;
  wire net_45554;
  wire net_45557;
  wire net_45560;
  wire net_45562;
  wire net_45563;
  wire net_45566;
  wire net_45568;
  wire net_45569;
  wire net_45570;
  wire net_45572;
  wire net_45574;
  wire net_45575;
  wire net_45576;
  wire net_45578;
  wire net_45580;
  wire net_45581;
  wire net_45582;
  wire net_45584;
  wire net_45586;
  wire net_45587;
  wire net_45588;
  wire net_45590;
  wire net_45592;
  wire net_45593;
  wire net_45594;
  wire net_45596;
  wire net_45598;
  wire net_45599;
  wire net_45600;
  wire net_45602;
  wire net_45604;
  wire net_45605;
  wire net_45606;
  wire net_45608;
  wire net_45609;
  wire net_45610;
  wire net_45612;
  wire net_45615;
  wire net_45616;
  wire net_45623;
  wire net_45627;
  wire net_45631;
  wire net_45632;
  wire net_45634;
  wire net_45646;
  wire net_45653;
  wire net_45654;
  wire net_45658;
  wire net_45662;
  wire net_45663;
  wire net_45665;
  wire net_45666;
  wire net_45683;
  wire net_45685;
  wire net_45687;
  wire net_45692;
  wire net_45693;
  wire net_45697;
  wire net_45702;
  wire net_45711;
  wire net_45715;
  wire net_45720;
  wire net_45727;
  wire net_45731;
  wire net_45732;
  wire net_45733;
  wire net_45734;
  wire net_45735;
  wire net_45736;
  wire net_45737;
  wire net_45738;
  wire net_45739;
  wire net_45740;
  wire net_45743;
  wire net_45747;
  wire net_45751;
  wire net_45757;
  wire net_45764;
  wire net_45767;
  wire net_45790;
  wire net_45791;
  wire net_45793;
  wire net_45796;
  wire net_45810;
  wire net_45814;
  wire net_45834;
  wire net_45850;
  wire net_45854;
  wire net_45855;
  wire net_45856;
  wire net_45857;
  wire net_45859;
  wire net_45860;
  wire net_45862;
  wire net_45863;
  wire net_45867;
  wire net_45872;
  wire net_45876;
  wire net_45879;
  wire net_45884;
  wire net_45885;
  wire net_45886;
  wire net_45888;
  wire net_45889;
  wire net_45905;
  wire net_45909;
  wire net_45923;
  wire net_45933;
  wire net_45957;
  wire net_45960;
  wire net_45976;
  wire net_45977;
  wire net_45979;
  wire net_45983;
  wire net_45984;
  wire net_45986;
  wire net_45988;
  wire net_45991;
  wire net_45993;
  wire net_45994;
  wire net_45996;
  wire net_46008;
  wire net_46011;
  wire net_46012;
  wire net_46021;
  wire net_46025;
  wire net_46028;
  wire net_46031;
  wire net_46033;
  wire net_46034;
  wire net_46040;
  wire net_46042;
  wire net_46043;
  wire net_46055;
  wire net_46061;
  wire net_46066;
  wire net_46071;
  wire net_46072;
  wire net_46079;
  wire net_46084;
  wire net_46086;
  wire net_46089;
  wire net_46092;
  wire net_46095;
  wire net_46096;
  wire net_46100;
  wire net_46101;
  wire net_46102;
  wire net_46107;
  wire net_46108;
  wire net_46114;
  wire net_46117;
  wire net_46119;
  wire net_46121;
  wire net_46124;
  wire net_46132;
  wire net_46136;
  wire net_46144;
  wire net_46154;
  wire net_46158;
  wire net_46183;
  wire net_46201;
  wire net_46221;
  wire net_46223;
  wire net_46224;
  wire net_46226;
  wire net_46228;
  wire net_46229;
  wire net_46231;
  wire net_46232;
  wire net_46235;
  wire net_46249;
  wire net_46250;
  wire net_46252;
  wire net_46258;
  wire net_46260;
  wire net_46268;
  wire net_46273;
  wire net_46283;
  wire net_46285;
  wire net_46307;
  wire net_46324;
  wire net_46343;
  wire net_46345;
  wire net_46346;
  wire net_46350;
  wire net_46351;
  wire net_46352;
  wire net_46353;
  wire net_46354;
  wire net_46358;
  wire net_46365;
  wire net_46369;
  wire net_46376;
  wire net_46389;
  wire net_46392;
  wire net_46395;
  wire net_46397;
  wire net_46401;
  wire net_46402;
  wire net_46403;
  wire net_46405;
  wire net_46409;
  wire net_46410;
  wire net_46414;
  wire net_46417;
  wire net_46422;
  wire net_46423;
  wire net_46424;
  wire net_46425;
  wire net_46429;
  wire net_46434;
  wire net_46437;
  wire net_46442;
  wire net_46443;
  wire net_46447;
  wire net_46455;
  wire net_46459;
  wire net_46465;
  wire net_46467;
  wire net_46469;
  wire net_46470;
  wire net_46471;
  wire net_46472;
  wire net_46474;
  wire net_46496;
  wire net_46503;
  wire net_46512;
  wire net_46518;
  wire net_46519;
  wire net_46522;
  wire net_46523;
  wire net_46527;
  wire net_46529;
  wire net_46530;
  wire net_46535;
  wire net_46536;
  wire net_46538;
  wire net_46540;
  wire net_46543;
  wire net_46546;
  wire net_46547;
  wire net_46548;
  wire net_46551;
  wire net_46552;
  wire net_46553;
  wire net_46557;
  wire net_46558;
  wire net_46560;
  wire net_46569;
  wire net_46570;
  wire net_46571;
  wire net_46572;
  wire net_46575;
  wire net_46576;
  wire net_46577;
  wire net_46591;
  wire net_46592;
  wire net_46593;
  wire net_46594;
  wire net_46596;
  wire net_46597;
  wire net_46598;
  wire net_46599;
  wire net_46600;
  wire net_46608;
  wire net_46610;
  wire net_46621;
  wire net_46627;
  wire net_46636;
  wire net_46644;
  wire net_46653;
  wire net_46655;
  wire net_46660;
  wire net_46661;
  wire net_46680;
  wire net_46681;
  wire net_46682;
  wire net_46683;
  wire net_46694;
  wire net_46714;
  wire net_46715;
  wire net_46717;
  wire net_46718;
  wire net_46720;
  wire net_46721;
  wire net_46722;
  wire net_46723;
  wire net_46730;
  wire net_46732;
  wire net_46740;
  wire net_46741;
  wire net_46743;
  wire net_46747;
  wire net_46749;
  wire net_46758;
  wire net_46761;
  wire net_46762;
  wire net_46768;
  wire net_46771;
  wire net_46785;
  wire net_46794;
  wire net_46806;
  wire net_46817;
  wire net_46824;
  wire net_46834;
  wire net_46837;
  wire net_46838;
  wire net_46840;
  wire net_46841;
  wire net_46842;
  wire net_46843;
  wire net_46844;
  wire net_46845;
  wire net_46847;
  wire net_46852;
  wire net_46854;
  wire net_46858;
  wire net_46875;
  wire net_46882;
  wire net_46885;
  wire net_46887;
  wire net_46896;
  wire net_46897;
  wire net_46899;
  wire net_46901;
  wire net_46902;
  wire net_46904;
  wire net_46910;
  wire net_46911;
  wire net_46915;
  wire net_46923;
  wire net_46926;
  wire net_46927;
  wire net_46928;
  wire net_46929;
  wire net_46938;
  wire net_46950;
  wire net_46956;
  wire net_46957;
  wire net_46958;
  wire net_46959;
  wire net_46960;
  wire net_46961;
  wire net_46963;
  wire net_46964;
  wire net_46965;
  wire net_46966;
  wire net_46967;
  wire net_46968;
  wire net_46969;
  wire net_46970;
  wire net_46976;
  wire net_46978;
  wire net_46986;
  wire net_46987;
  wire net_46989;
  wire net_46997;
  wire net_47008;
  wire net_47012;
  wire net_47013;
  wire net_47018;
  wire net_47022;
  wire net_47023;
  wire net_47030;
  wire net_47031;
  wire net_47033;
  wire net_47037;
  wire net_47038;
  wire net_47039;
  wire net_47043;
  wire net_47045;
  wire net_47046;
  wire net_47055;
  wire net_47056;
  wire net_47057;
  wire net_47062;
  wire net_47063;
  wire net_47064;
  wire net_47083;
  wire net_47084;
  wire net_47085;
  wire net_47087;
  wire net_47088;
  wire net_47089;
  wire net_47090;
  wire net_47092;
  wire net_47093;
  wire net_47113;
  wire net_47119;
  wire net_47128;
  wire net_47129;
  wire net_47131;
  wire net_47132;
  wire net_47135;
  wire net_47136;
  wire net_47137;
  wire net_47138;
  wire net_47141;
  wire net_47143;
  wire net_47145;
  wire net_47156;
  wire net_47162;
  wire net_47173;
  wire net_47181;
  wire net_47185;
  wire net_47190;
  wire net_47191;
  wire net_47192;
  wire net_47193;
  wire net_47196;
  wire net_47197;
  wire net_47198;
  wire net_47199;
  wire net_47205;
  wire net_47206;
  wire net_47207;
  wire net_47211;
  wire net_47213;
  wire net_47229;
  wire net_47235;
  wire net_47250;
  wire net_47251;
  wire net_47252;
  wire net_47255;
  wire net_47256;
  wire net_47257;
  wire net_47260;
  wire net_47263;
  wire net_47264;
  wire net_47265;
  wire net_47266;
  wire net_47268;
  wire net_47277;
  wire net_47278;
  wire net_47280;
  wire net_47289;
  wire net_47290;
  wire net_47291;
  wire net_47292;
  wire net_47295;
  wire net_47296;
  wire net_47297;
  wire net_47298;
  wire net_47313;
  wire net_47314;
  wire net_47315;
  wire net_47316;
  wire net_47325;
  wire net_47326;
  wire net_47327;
  wire net_47328;
  wire net_47329;
  wire net_47330;
  wire net_47335;
  wire net_47382;
  wire net_47413;
  wire net_47452;
  wire net_47453;
  wire net_48810;
  wire net_48880;
  wire net_48911;
  wire net_48913;
  wire net_48914;
  wire net_48926;
  wire net_48932;
  wire net_48952;
  wire net_48954;
  wire net_48959;
  wire net_48967;
  wire net_48968;
  wire net_48975;
  wire net_48977;
  wire net_48979;
  wire net_48985;
  wire net_48988;
  wire net_48989;
  wire net_48990;
  wire net_48992;
  wire net_48994;
  wire net_48995;
  wire net_48997;
  wire net_48998;
  wire net_49000;
  wire net_49001;
  wire net_49002;
  wire net_49004;
  wire net_49008;
  wire net_49009;
  wire net_49010;
  wire net_49029;
  wire net_49030;
  wire net_49031;
  wire net_49034;
  wire net_49036;
  wire net_49037;
  wire net_49038;
  wire net_49039;
  wire net_49040;
  wire net_49051;
  wire net_49071;
  wire net_49073;
  wire net_49074;
  wire net_49076;
  wire net_49078;
  wire net_49089;
  wire net_49090;
  wire net_49091;
  wire net_49092;
  wire net_49093;
  wire net_49094;
  wire net_49096;
  wire net_49115;
  wire net_49119;
  wire net_49123;
  wire net_49124;
  wire net_49131;
  wire net_49134;
  wire net_49148;
  wire net_49155;
  wire net_49158;
  wire net_49164;
  wire net_49170;
  wire net_49183;
  wire net_49193;
  wire net_49194;
  wire net_49195;
  wire net_49196;
  wire net_49197;
  wire net_49199;
  wire net_49200;
  wire net_49201;
  wire net_49202;
  wire net_49211;
  wire net_49219;
  wire net_49224;
  wire net_49230;
  wire net_49236;
  wire net_49238;
  wire net_49239;
  wire net_49240;
  wire net_49241;
  wire net_49246;
  wire net_49256;
  wire net_49257;
  wire net_49258;
  wire net_49266;
  wire net_49271;
  wire net_49276;
  wire net_49282;
  wire net_49286;
  wire net_49289;
  wire net_49294;
  wire net_49295;
  wire net_49296;
  wire net_49299;
  wire net_49308;
  wire net_49312;
  wire net_49314;
  wire net_49316;
  wire net_49317;
  wire net_49318;
  wire net_49319;
  wire net_49320;
  wire net_49321;
  wire net_49322;
  wire net_49323;
  wire net_49324;
  wire net_49325;
  wire net_49337;
  wire net_49340;
  wire net_49343;
  wire net_49346;
  wire net_49351;
  wire net_49363;
  wire net_49365;
  wire net_49366;
  wire net_49367;
  wire net_49371;
  wire net_49373;
  wire net_49375;
  wire net_49378;
  wire net_49379;
  wire net_49380;
  wire net_49383;
  wire net_49384;
  wire net_49385;
  wire net_49386;
  wire net_49388;
  wire net_49390;
  wire net_49395;
  wire net_49398;
  wire net_49399;
  wire net_49400;
  wire net_49401;
  wire net_49405;
  wire net_49410;
  wire net_49418;
  wire net_49422;
  wire net_49425;
  wire net_49428;
  wire net_49429;
  wire net_49430;
  wire net_49431;
  wire net_49435;
  wire net_49437;
  wire net_49438;
  wire net_49439;
  wire net_49441;
  wire net_49442;
  wire net_49446;
  wire net_49447;
  wire net_49456;
  wire net_49460;
  wire net_49461;
  wire net_49464;
  wire net_49467;
  wire net_49468;
  wire net_49469;
  wire net_49493;
  wire net_49494;
  wire net_49495;
  wire net_49511;
  wire net_49517;
  wire net_49527;
  wire net_49546;
  wire net_49552;
  wire net_49561;
  wire net_49562;
  wire net_49564;
  wire net_49565;
  wire net_49566;
  wire net_49567;
  wire net_49568;
  wire net_49569;
  wire net_49570;
  wire net_49571;
  wire net_49576;
  wire net_49578;
  wire net_49608;
  wire net_49610;
  wire net_49616;
  wire net_49617;
  wire net_49620;
  wire net_49623;
  wire net_49629;
  wire net_49630;
  wire net_49636;
  wire net_49640;
  wire net_49645;
  wire net_49653;
  wire net_49656;
  wire net_49663;
  wire net_49665;
  wire net_49670;
  wire net_49671;
  wire net_49674;
  wire net_49677;
  wire net_49683;
  wire net_49685;
  wire net_49686;
  wire net_49687;
  wire net_49688;
  wire net_49689;
  wire net_49690;
  wire net_49691;
  wire net_49692;
  wire net_49693;
  wire net_49694;
  wire net_49698;
  wire net_49704;
  wire net_49708;
  wire net_49710;
  wire net_49737;
  wire net_49739;
  wire net_49741;
  wire net_49742;
  wire net_49744;
  wire net_49745;
  wire net_49750;
  wire net_49752;
  wire net_49755;
  wire net_49763;
  wire net_49767;
  wire net_49779;
  wire net_49780;
  wire net_49781;
  wire net_49782;
  wire net_49785;
  wire net_49797;
  wire net_49804;
  wire net_49807;
  wire net_49808;
  wire net_49810;
  wire net_49811;
  wire net_49812;
  wire net_49814;
  wire net_49815;
  wire net_49816;
  wire net_49817;
  wire net_49827;
  wire net_49828;
  wire net_49836;
  wire net_49841;
  wire net_49855;
  wire net_49857;
  wire net_49859;
  wire net_49861;
  wire net_49886;
  wire net_49909;
  wire net_49916;
  wire net_49927;
  wire net_49930;
  wire net_49931;
  wire net_49935;
  wire net_49938;
  wire net_49945;
  wire net_49952;
  wire net_49955;
  wire net_49956;
  wire net_49968;
  wire net_49985;
  wire net_49993;
  wire net_49998;
  wire net_50001;
  wire net_50010;
  wire net_50038;
  wire net_50046;
  wire net_50053;
  wire net_50054;
  wire net_50056;
  wire net_50057;
  wire net_50058;
  wire net_50060;
  wire net_50061;
  wire net_50086;
  wire net_50087;
  wire net_50091;
  wire net_50097;
  wire net_50100;
  wire net_50101;
  wire net_50108;
  wire net_50110;
  wire net_50122;
  wire net_50139;
  wire net_50149;
  wire net_50151;
  wire net_50154;
  wire net_50166;
  wire net_50168;
  wire net_50174;
  wire net_50177;
  wire net_50178;
  wire net_50180;
  wire net_50181;
  wire net_50183;
  wire net_50184;
  wire net_50185;
  wire net_50206;
  wire net_50207;
  wire net_50212;
  wire net_50214;
  wire net_50222;
  wire net_50224;
  wire net_50227;
  wire net_50231;
  wire net_50233;
  wire net_50235;
  wire net_50265;
  wire net_50274;
  wire net_50279;
  wire net_50285;
  wire net_50291;
  wire net_50299;
  wire net_50300;
  wire net_50302;
  wire net_50303;
  wire net_50304;
  wire net_50305;
  wire net_50306;
  wire net_50307;
  wire net_50308;
  wire net_50309;
  wire net_50314;
  wire net_50320;
  wire net_50323;
  wire net_50327;
  wire net_50331;
  wire net_50333;
  wire net_50334;
  wire net_50335;
  wire net_50345;
  wire net_50353;
  wire net_50355;
  wire net_50362;
  wire net_50363;
  wire net_50368;
  wire net_50372;
  wire net_50379;
  wire net_50383;
  wire net_50394;
  wire net_50395;
  wire net_50396;
  wire net_50397;
  wire net_50422;
  wire net_50423;
  wire net_50425;
  wire net_50426;
  wire net_50427;
  wire net_50428;
  wire net_50429;
  wire net_50430;
  wire net_50431;
  wire net_50432;
  wire net_50445;
  wire net_50450;
  wire net_50451;
  wire net_50453;
  wire net_50455;
  wire net_50460;
  wire net_50466;
  wire net_50472;
  wire net_50475;
  wire net_50476;
  wire net_50477;
  wire net_50492;
  wire net_50494;
  wire net_50501;
  wire net_50514;
  wire net_50517;
  wire net_50518;
  wire net_50523;
  wire net_50532;
  wire net_50538;
  wire net_50546;
  wire net_50547;
  wire net_50548;
  wire net_50549;
  wire net_50550;
  wire net_50551;
  wire net_50552;
  wire net_50553;
  wire net_50554;
  wire net_50555;
  wire net_50567;
  wire net_50573;
  wire net_50575;
  wire net_50578;
  wire net_50579;
  wire net_50580;
  wire net_50581;
  wire net_50583;
  wire net_50590;
  wire net_50598;
  wire net_50599;
  wire net_50600;
  wire net_50602;
  wire net_50606;
  wire net_50609;
  wire net_50612;
  wire net_50614;
  wire net_50616;
  wire net_50617;
  wire net_50619;
  wire net_50622;
  wire net_50624;
  wire net_50625;
  wire net_50628;
  wire net_50629;
  wire net_50630;
  wire net_50640;
  wire net_50642;
  wire net_50643;
  wire net_50647;
  wire net_50648;
  wire net_50649;
  wire net_50652;
  wire net_50654;
  wire net_50658;
  wire net_50659;
  wire net_50661;
  wire net_50668;
  wire net_50669;
  wire net_50670;
  wire net_50671;
  wire net_50672;
  wire net_50673;
  wire net_50675;
  wire net_50676;
  wire net_50677;
  wire net_50678;
  wire net_50686;
  wire net_50691;
  wire net_50692;
  wire net_50697;
  wire net_50701;
  wire net_50714;
  wire net_50715;
  wire net_50723;
  wire net_50724;
  wire net_50731;
  wire net_50734;
  wire net_50739;
  wire net_50740;
  wire net_50742;
  wire net_50748;
  wire net_50751;
  wire net_50752;
  wire net_50753;
  wire net_50754;
  wire net_50757;
  wire net_50758;
  wire net_50759;
  wire net_50760;
  wire net_50763;
  wire net_50764;
  wire net_50765;
  wire net_50766;
  wire net_50770;
  wire net_50771;
  wire net_50772;
  wire net_50775;
  wire net_50776;
  wire net_50777;
  wire net_50787;
  wire net_50788;
  wire net_50789;
  wire net_50790;
  wire net_50791;
  wire net_50792;
  wire net_50793;
  wire net_50795;
  wire net_50796;
  wire net_50797;
  wire net_50798;
  wire net_50799;
  wire net_50800;
  wire net_50801;
  wire net_50806;
  wire net_50812;
  wire net_50820;
  wire net_50821;
  wire net_50828;
  wire net_50835;
  wire net_50836;
  wire net_50837;
  wire net_50838;
  wire net_50839;
  wire net_50840;
  wire net_50841;
  wire net_50842;
  wire net_50844;
  wire net_50846;
  wire net_50847;
  wire net_50848;
  wire net_50849;
  wire net_50850;
  wire net_50856;
  wire net_50857;
  wire net_50858;
  wire net_50864;
  wire net_50866;
  wire net_50868;
  wire net_50869;
  wire net_50870;
  wire net_50871;
  wire net_50874;
  wire net_50875;
  wire net_50876;
  wire net_50877;
  wire net_50880;
  wire net_50882;
  wire net_50886;
  wire net_50887;
  wire net_50888;
  wire net_50889;
  wire net_50894;
  wire net_50898;
  wire net_50899;
  wire net_50900;
  wire net_50901;
  wire net_50904;
  wire net_50905;
  wire net_50906;
  wire net_50907;
  wire net_50910;
  wire net_50911;
  wire net_50912;
  wire net_50913;
  wire net_50915;
  wire net_50916;
  wire net_50918;
  wire net_50920;
  wire net_50921;
  wire net_50922;
  wire net_50924;
  wire net_50929;
  wire net_50932;
  wire net_50943;
  wire net_50948;
  wire net_50959;
  wire net_50966;
  wire net_50971;
  wire net_50978;
  wire net_50993;
  wire net_50996;
  wire net_50999;
  wire net_51000;
  wire net_51003;
  wire net_51006;
  wire net_51011;
  wire net_51016;
  wire net_51027;
  wire net_51035;
  wire net_51038;
  wire net_51039;
  wire net_51040;
  wire net_51041;
  wire net_51042;
  wire net_51043;
  wire net_51045;
  wire net_51046;
  wire net_51047;
  wire net_51057;
  wire net_51066;
  wire net_51067;
  wire net_51073;
  wire net_51082;
  wire net_51092;
  wire net_51093;
  wire net_51129;
  wire net_51139;
  wire net_51160;
  wire net_51161;
  wire net_51170;
  wire net_51180;
  wire net_51218;
  wire net_51231;
  wire net_51255;
  wire net_51283;
  wire net_51284;
  wire net_52745;
  wire net_52762;
  wire net_52784;
  wire net_52785;
  wire net_52791;
  wire net_52792;
  wire net_52793;
  wire net_52832;
  wire net_52846;
  wire net_52847;
  wire net_52850;
  wire net_52851;
  wire net_52852;
  wire net_52861;
  wire net_52862;
  wire net_52867;
  wire net_52869;
  wire net_52870;
  wire net_52873;
  wire net_52921;
  wire net_52948;
  wire net_52952;
  wire net_52954;
  wire net_52955;
  wire net_52959;
  wire net_52963;
  wire net_52970;
  wire net_52971;
  wire net_52977;
  wire net_52980;
  wire net_52984;
  wire net_52985;
  wire net_52986;
  wire net_52990;
  wire net_52995;
  wire net_52998;
  wire net_53002;
  wire net_53023;
  wire net_53024;
  wire net_53025;
  wire net_53032;
  wire net_53033;
  wire net_53051;
  wire net_53053;
  wire net_53060;
  wire net_53067;
  wire net_53068;
  wire net_53070;
  wire net_53073;
  wire net_53074;
  wire net_53080;
  wire net_53083;
  wire net_53087;
  wire net_53088;
  wire net_53092;
  wire net_53093;
  wire net_53101;
  wire net_53109;
  wire net_53112;
  wire net_53126;
  wire net_53127;
  wire net_53131;
  wire net_53132;
  wire net_53138;
  wire net_53142;
  wire net_53144;
  wire net_53145;
  wire net_53147;
  wire net_53148;
  wire net_53149;
  wire net_53151;
  wire net_53152;
  wire net_53153;
  wire net_53154;
  wire net_53155;
  wire net_53156;
  wire net_53162;
  wire net_53163;
  wire net_53165;
  wire net_53179;
  wire net_53183;
  wire net_53192;
  wire net_53193;
  wire net_53194;
  wire net_53195;
  wire net_53198;
  wire net_53199;
  wire net_53200;
  wire net_53201;
  wire net_53203;
  wire net_53206;
  wire net_53207;
  wire net_53210;
  wire net_53211;
  wire net_53217;
  wire net_53223;
  wire net_53231;
  wire net_53235;
  wire net_53241;
  wire net_53242;
  wire net_53244;
  wire net_53248;
  wire net_53256;
  wire net_53259;
  wire net_53260;
  wire net_53261;
  wire net_53262;
  wire net_53265;
  wire net_53268;
  wire net_53270;
  wire net_53271;
  wire net_53272;
  wire net_53273;
  wire net_53274;
  wire net_53275;
  wire net_53276;
  wire net_53277;
  wire net_53278;
  wire net_53279;
  wire net_53284;
  wire net_53286;
  wire net_53288;
  wire net_53290;
  wire net_53294;
  wire net_53295;
  wire net_53296;
  wire net_53301;
  wire net_53315;
  wire net_53322;
  wire net_53324;
  wire net_53331;
  wire net_53332;
  wire net_53346;
  wire net_53354;
  wire net_53377;
  wire net_53384;
  wire net_53392;
  wire net_53393;
  wire net_53395;
  wire net_53396;
  wire net_53398;
  wire net_53399;
  wire net_53400;
  wire net_53401;
  wire net_53402;
  wire net_53407;
  wire net_53411;
  wire net_53415;
  wire net_53428;
  wire net_53439;
  wire net_53441;
  wire net_53445;
  wire net_53450;
  wire net_53451;
  wire net_53453;
  wire net_53454;
  wire net_53455;
  wire net_53458;
  wire net_53462;
  wire net_53467;
  wire net_53472;
  wire net_53475;
  wire net_53484;
  wire net_53487;
  wire net_53493;
  wire net_53494;
  wire net_53495;
  wire net_53496;
  wire net_53500;
  wire net_53505;
  wire net_53512;
  wire net_53515;
  wire net_53516;
  wire net_53519;
  wire net_53521;
  wire net_53523;
  wire net_53524;
  wire net_53525;
  wire net_53529;
  wire net_53530;
  wire net_53532;
  wire net_53534;
  wire net_53540;
  wire net_53550;
  wire net_53552;
  wire net_53559;
  wire net_53564;
  wire net_53566;
  wire net_53567;
  wire net_53569;
  wire net_53570;
  wire net_53578;
  wire net_53579;
  wire net_53580;
  wire net_53584;
  wire net_53586;
  wire net_53587;
  wire net_53588;
  wire net_53589;
  wire net_53590;
  wire net_53595;
  wire net_53600;
  wire net_53604;
  wire net_53605;
  wire net_53606;
  wire net_53607;
  wire net_53610;
  wire net_53616;
  wire net_53624;
  wire net_53630;
  wire net_53634;
  wire net_53635;
  wire net_53636;
  wire net_53637;
  wire net_53638;
  wire net_53639;
  wire net_53641;
  wire net_53642;
  wire net_53643;
  wire net_53644;
  wire net_53645;
  wire net_53646;
  wire net_53647;
  wire net_53648;
  wire net_53651;
  wire net_53654;
  wire net_53657;
  wire net_53666;
  wire net_53670;
  wire net_53672;
  wire net_53673;
  wire net_53674;
  wire net_53682;
  wire net_53684;
  wire net_53685;
  wire net_53686;
  wire net_53687;
  wire net_53688;
  wire net_53691;
  wire net_53692;
  wire net_53693;
  wire net_53695;
  wire net_53696;
  wire net_53699;
  wire net_53701;
  wire net_53702;
  wire net_53703;
  wire net_53711;
  wire net_53712;
  wire net_53715;
  wire net_53716;
  wire net_53717;
  wire net_53718;
  wire net_53721;
  wire net_53722;
  wire net_53723;
  wire net_53724;
  wire net_53727;
  wire net_53728;
  wire net_53729;
  wire net_53739;
  wire net_53741;
  wire net_53742;
  wire net_53745;
  wire net_53746;
  wire net_53747;
  wire net_53751;
  wire net_53753;
  wire net_53754;
  wire net_53757;
  wire net_53758;
  wire net_53760;
  wire net_53761;
  wire net_53762;
  wire net_53763;
  wire net_53764;
  wire net_53765;
  wire net_53770;
  wire net_53774;
  wire net_53776;
  wire net_53777;
  wire net_53778;
  wire net_53779;
  wire net_53780;
  wire net_53788;
  wire net_53798;
  wire net_53811;
  wire net_53816;
  wire net_53832;
  wire net_53852;
  wire net_53871;
  wire net_53884;
  wire net_53885;
  wire net_53887;
  wire net_53888;
  wire net_53889;
  wire net_53890;
  wire net_53891;
  wire net_53892;
  wire net_53893;
  wire net_53894;
  wire net_53897;
  wire net_53898;
  wire net_53902;
  wire net_53905;
  wire net_53908;
  wire net_53909;
  wire net_53911;
  wire net_53920;
  wire net_53929;
  wire net_53940;
  wire net_53941;
  wire net_53942;
  wire net_53944;
  wire net_53945;
  wire net_53946;
  wire net_53949;
  wire net_53952;
  wire net_53953;
  wire net_53955;
  wire net_53961;
  wire net_53962;
  wire net_53963;
  wire net_53964;
  wire net_53969;
  wire net_53974;
  wire net_53985;
  wire net_53986;
  wire net_53987;
  wire net_53988;
  wire net_53991;
  wire net_54007;
  wire net_54008;
  wire net_54010;
  wire net_54013;
  wire net_54014;
  wire net_54017;
  wire net_54019;
  wire net_54025;
  wire net_54027;
  wire net_54029;
  wire net_54030;
  wire net_54031;
  wire net_54033;
  wire net_54055;
  wire net_54056;
  wire net_54058;
  wire net_54066;
  wire net_54070;
  wire net_54072;
  wire net_54073;
  wire net_54078;
  wire net_54082;
  wire net_54093;
  wire net_54099;
  wire net_54108;
  wire net_54109;
  wire net_54110;
  wire net_54111;
  wire net_54116;
  wire net_54122;
  wire net_54130;
  wire net_54131;
  wire net_54137;
  wire net_54144;
  wire net_54146;
  wire net_54151;
  wire net_54155;
  wire net_54159;
  wire net_54163;
  wire net_54176;
  wire net_54179;
  wire net_54180;
  wire net_54183;
  wire net_54184;
  wire net_54195;
  wire net_54196;
  wire net_54199;
  wire net_54205;
  wire net_54207;
  wire net_54216;
  wire net_54220;
  wire net_54228;
  wire net_54232;
  wire net_54240;
  wire net_54245;
  wire net_54251;
  wire net_54253;
  wire net_54254;
  wire net_54256;
  wire net_54257;
  wire net_54258;
  wire net_54259;
  wire net_54260;
  wire net_54261;
  wire net_54262;
  wire net_54263;
  wire net_54284;
  wire net_54286;
  wire net_54289;
  wire net_54299;
  wire net_54303;
  wire net_54304;
  wire net_54305;
  wire net_54307;
  wire net_54308;
  wire net_54309;
  wire net_54311;
  wire net_54313;
  wire net_54316;
  wire net_54317;
  wire net_54323;
  wire net_54324;
  wire net_54325;
  wire net_54326;
  wire net_54331;
  wire net_54336;
  wire net_54337;
  wire net_54338;
  wire net_54339;
  wire net_54345;
  wire net_54351;
  wire net_54354;
  wire net_54355;
  wire net_54356;
  wire net_54357;
  wire net_54360;
  wire net_54366;
  wire net_54367;
  wire net_54368;
  wire net_54369;
  wire net_54372;
  wire net_54373;
  wire net_54374;
  wire net_54375;
  wire net_54376;
  wire net_54377;
  wire net_54379;
  wire net_54381;
  wire net_54383;
  wire net_54384;
  wire net_54385;
  wire net_54386;
  wire net_54396;
  wire net_54408;
  wire net_54409;
  wire net_54411;
  wire net_54413;
  wire net_54425;
  wire net_54427;
  wire net_54428;
  wire net_54429;
  wire net_54431;
  wire net_54433;
  wire net_54435;
  wire net_54436;
  wire net_54437;
  wire net_54438;
  wire net_54444;
  wire net_54446;
  wire net_54447;
  wire net_54450;
  wire net_54453;
  wire net_54459;
  wire net_54461;
  wire net_54465;
  wire net_54466;
  wire net_54471;
  wire net_54478;
  wire net_54486;
  wire net_54491;
  wire net_54495;
  wire net_54496;
  wire net_54497;
  wire net_54498;
  wire net_54499;
  wire net_54500;
  wire net_54502;
  wire net_54503;
  wire net_54504;
  wire net_54505;
  wire net_54506;
  wire net_54507;
  wire net_54508;
  wire net_54509;
  wire net_54514;
  wire net_54516;
  wire net_54518;
  wire net_54520;
  wire net_54543;
  wire net_54544;
  wire net_54546;
  wire net_54549;
  wire net_54551;
  wire net_54552;
  wire net_54553;
  wire net_54554;
  wire net_54555;
  wire net_54556;
  wire net_54561;
  wire net_54567;
  wire net_54574;
  wire net_54576;
  wire net_54578;
  wire net_54582;
  wire net_54584;
  wire net_54585;
  wire net_54588;
  wire net_54589;
  wire net_54590;
  wire net_54591;
  wire net_54603;
  wire net_54607;
  wire net_54615;
  wire net_54620;
  wire net_54622;
  wire net_54623;
  wire net_54627;
  wire net_54628;
  wire net_54629;
  wire net_54630;
  wire net_54631;
  wire net_54632;
  wire net_54652;
  wire net_54654;
  wire net_54656;
  wire net_54658;
  wire net_54660;
  wire net_54667;
  wire net_54668;
  wire net_54669;
  wire net_54670;
  wire net_54672;
  wire net_54673;
  wire net_54676;
  wire net_54677;
  wire net_54678;
  wire net_54679;
  wire net_54682;
  wire net_54685;
  wire net_54694;
  wire net_54695;
  wire net_54696;
  wire net_54700;
  wire net_54704;
  wire net_54707;
  wire net_54708;
  wire net_54711;
  wire net_54714;
  wire net_54719;
  wire net_54720;
  wire net_54723;
  wire net_54724;
  wire net_54725;
  wire net_54726;
  wire net_54729;
  wire net_54730;
  wire net_54731;
  wire net_54735;
  wire net_54736;
  wire net_54737;
  wire net_54738;
  wire net_54742;
  wire net_54746;
  wire net_54747;
  wire net_54748;
  wire net_54749;
  wire net_54750;
  wire net_54751;
  wire net_54753;
  wire net_54754;
  wire net_54755;
  wire net_54765;
  wire net_54771;
  wire net_54772;
  wire net_54775;
  wire net_54780;
  wire net_54789;
  wire net_54790;
  wire net_54793;
  wire net_54796;
  wire net_54800;
  wire net_54803;
  wire net_54804;
  wire net_54816;
  wire net_54828;
  wire net_54829;
  wire net_54831;
  wire net_54842;
  wire net_54847;
  wire net_54852;
  wire net_54853;
  wire net_54854;
  wire net_54855;
  wire net_54865;
  wire net_54869;
  wire net_54870;
  wire net_54871;
  wire net_54872;
  wire net_54873;
  wire net_54874;
  wire net_54876;
  wire net_54877;
  wire net_54878;
  wire net_54888;
  wire net_54905;
  wire net_54912;
  wire net_54913;
  wire net_54915;
  wire net_54916;
  wire net_54917;
  wire net_54919;
  wire net_54920;
  wire net_54923;
  wire net_54924;
  wire net_54925;
  wire net_54926;
  wire net_54927;
  wire net_54928;
  wire net_54929;
  wire net_54930;
  wire net_54931;
  wire net_54933;
  wire net_54935;
  wire net_54936;
  wire net_54938;
  wire net_54939;
  wire net_54941;
  wire net_54942;
  wire net_54945;
  wire net_54946;
  wire net_54947;
  wire net_54948;
  wire net_54951;
  wire net_54952;
  wire net_54953;
  wire net_54954;
  wire net_54957;
  wire net_54958;
  wire net_54959;
  wire net_54960;
  wire net_54963;
  wire net_54964;
  wire net_54965;
  wire net_54966;
  wire net_54975;
  wire net_54976;
  wire net_54977;
  wire net_54978;
  wire net_54981;
  wire net_54982;
  wire net_54983;
  wire net_54984;
  wire net_54987;
  wire net_54988;
  wire net_54989;
  wire net_54990;
  wire net_54991;
  wire net_54992;
  wire net_54997;
  wire net_55036;
  wire net_55039;
  wire net_55044;
  wire net_55046;
  wire net_55049;
  wire net_55110;
  wire net_55111;
  wire net_55112;
  wire net_55113;
  wire net_55114;
  wire net_55115;
  wire net_56515;
  wire net_56518;
  wire net_56527;
  wire net_56533;
  wire net_56601;
  wire net_56614;
  wire net_56627;
  wire net_56682;
  wire net_56683;
  wire net_56693;
  wire net_56703;
  wire net_56738;
  wire net_56757;
  wire net_56774;
  wire net_56776;
  wire net_56779;
  wire net_56783;
  wire net_56785;
  wire net_56788;
  wire net_56809;
  wire net_56820;
  wire net_56826;
  wire net_56827;
  wire net_56828;
  wire net_56845;
  wire net_56853;
  wire net_56854;
  wire net_56855;
  wire net_56858;
  wire net_56860;
  wire net_56883;
  wire net_56889;
  wire net_56900;
  wire net_56907;
  wire net_56969;
  wire net_56972;
  wire net_56976;
  wire net_56977;
  wire net_56978;
  wire net_56979;
  wire net_56980;
  wire net_56981;
  wire net_56982;
  wire net_56983;
  wire net_56984;
  wire net_56985;
  wire net_56986;
  wire net_56992;
  wire net_57003;
  wire net_57007;
  wire net_57008;
  wire net_57009;
  wire net_57020;
  wire net_57026;
  wire net_57032;
  wire net_57035;
  wire net_57040;
  wire net_57043;
  wire net_57045;
  wire net_57048;
  wire net_57051;
  wire net_57055;
  wire net_57065;
  wire net_57066;
  wire net_57067;
  wire net_57071;
  wire net_57079;
  wire net_57083;
  wire net_57089;
  wire net_57096;
  wire net_57099;
  wire net_57100;
  wire net_57102;
  wire net_57103;
  wire net_57104;
  wire net_57105;
  wire net_57106;
  wire net_57107;
  wire net_57108;
  wire net_57109;
  wire net_57126;
  wire net_57134;
  wire net_57135;
  wire net_57137;
  wire net_57143;
  wire net_57145;
  wire net_57146;
  wire net_57152;
  wire net_57155;
  wire net_57156;
  wire net_57159;
  wire net_57160;
  wire net_57162;
  wire net_57163;
  wire net_57165;
  wire net_57166;
  wire net_57168;
  wire net_57170;
  wire net_57172;
  wire net_57173;
  wire net_57174;
  wire net_57176;
  wire net_57177;
  wire net_57178;
  wire net_57179;
  wire net_57183;
  wire net_57188;
  wire net_57197;
  wire net_57200;
  wire net_57201;
  wire net_57202;
  wire net_57203;
  wire net_57206;
  wire net_57207;
  wire net_57208;
  wire net_57209;
  wire net_57214;
  wire net_57218;
  wire net_57222;
  wire net_57223;
  wire net_57225;
  wire net_57226;
  wire net_57228;
  wire net_57229;
  wire net_57230;
  wire net_57231;
  wire net_57232;
  wire net_57250;
  wire net_57266;
  wire net_57269;
  wire net_57270;
  wire net_57273;
  wire net_57275;
  wire net_57276;
  wire net_57277;
  wire net_57278;
  wire net_57279;
  wire net_57282;
  wire net_57288;
  wire net_57290;
  wire net_57294;
  wire net_57295;
  wire net_57296;
  wire net_57302;
  wire net_57305;
  wire net_57306;
  wire net_57307;
  wire net_57308;
  wire net_57317;
  wire net_57318;
  wire net_57319;
  wire net_57320;
  wire net_57325;
  wire net_57326;
  wire net_57332;
  wire net_57337;
  wire net_57341;
  wire net_57342;
  wire net_57343;
  wire net_57344;
  wire net_57346;
  wire net_57347;
  wire net_57350;
  wire net_57351;
  wire net_57352;
  wire net_57354;
  wire net_57356;
  wire net_57360;
  wire net_57364;
  wire net_57366;
  wire net_57370;
  wire net_57396;
  wire net_57402;
  wire net_57404;
  wire net_57407;
  wire net_57416;
  wire net_57429;
  wire net_57440;
  wire net_57455;
  wire net_57460;
  wire net_57465;
  wire net_57469;
  wire net_57470;
  wire net_57471;
  wire net_57472;
  wire net_57473;
  wire net_57474;
  wire net_57475;
  wire net_57482;
  wire net_57486;
  wire net_57491;
  wire net_57504;
  wire net_57512;
  wire net_57513;
  wire net_57517;
  wire net_57521;
  wire net_57523;
  wire net_57524;
  wire net_57525;
  wire net_57528;
  wire net_57536;
  wire net_57538;
  wire net_57541;
  wire net_57547;
  wire net_57552;
  wire net_57559;
  wire net_57563;
  wire net_57570;
  wire net_57576;
  wire net_57581;
  wire net_57582;
  wire net_57583;
  wire net_57584;
  wire net_57587;
  wire net_57592;
  wire net_57593;
  wire net_57594;
  wire net_57595;
  wire net_57596;
  wire net_57597;
  wire net_57598;
  wire net_57600;
  wire net_57603;
  wire net_57605;
  wire net_57606;
  wire net_57607;
  wire net_57609;
  wire net_57610;
  wire net_57613;
  wire net_57617;
  wire net_57618;
  wire net_57619;
  wire net_57621;
  wire net_57629;
  wire net_57635;
  wire net_57636;
  wire net_57637;
  wire net_57639;
  wire net_57643;
  wire net_57644;
  wire net_57646;
  wire net_57668;
  wire net_57675;
  wire net_57704;
  wire net_57705;
  wire net_57706;
  wire net_57707;
  wire net_57714;
  wire net_57715;
  wire net_57718;
  wire net_57719;
  wire net_57720;
  wire net_57723;
  wire net_57724;
  wire net_57729;
  wire net_57731;
  wire net_57741;
  wire net_57743;
  wire net_57744;
  wire net_57745;
  wire net_57746;
  wire net_57747;
  wire net_57750;
  wire net_57751;
  wire net_57752;
  wire net_57759;
  wire net_57760;
  wire net_57771;
  wire net_57773;
  wire net_57774;
  wire net_57778;
  wire net_57781;
  wire net_57782;
  wire net_57786;
  wire net_57792;
  wire net_57794;
  wire net_57797;
  wire net_57799;
  wire net_57803;
  wire net_57804;
  wire net_57809;
  wire net_57810;
  wire net_57817;
  wire net_57821;
  wire net_57824;
  wire net_57828;
  wire net_57830;
  wire net_57834;
  wire net_57835;
  wire net_57838;
  wire net_57839;
  wire net_57840;
  wire net_57841;
  wire net_57842;
  wire net_57843;
  wire net_57844;
  wire net_57845;
  wire net_57846;
  wire net_57847;
  wire net_57883;
  wire net_57884;
  wire net_57890;
  wire net_57893;
  wire net_57896;
  wire net_57914;
  wire net_57934;
  wire net_57939;
  wire net_57959;
  wire net_57960;
  wire net_57961;
  wire net_57963;
  wire net_57964;
  wire net_57965;
  wire net_57966;
  wire net_57967;
  wire net_57968;
  wire net_57969;
  wire net_57970;
  wire net_57975;
  wire net_57978;
  wire net_57982;
  wire net_57987;
  wire net_57990;
  wire net_57995;
  wire net_57996;
  wire net_57998;
  wire net_58012;
  wire net_58062;
  wire net_58084;
  wire net_58085;
  wire net_58087;
  wire net_58088;
  wire net_58089;
  wire net_58090;
  wire net_58091;
  wire net_58092;
  wire net_58093;
  wire net_58096;
  wire net_58106;
  wire net_58110;
  wire net_58114;
  wire net_58115;
  wire net_58116;
  wire net_58131;
  wire net_58133;
  wire net_58139;
  wire net_58143;
  wire net_58144;
  wire net_58145;
  wire net_58147;
  wire net_58151;
  wire net_58152;
  wire net_58154;
  wire net_58155;
  wire net_58160;
  wire net_58167;
  wire net_58174;
  wire net_58178;
  wire net_58179;
  wire net_58180;
  wire net_58186;
  wire net_58193;
  wire net_58196;
  wire net_58197;
  wire net_58198;
  wire net_58199;
  wire net_58204;
  wire net_58207;
  wire net_58208;
  wire net_58209;
  wire net_58210;
  wire net_58211;
  wire net_58212;
  wire net_58213;
  wire net_58214;
  wire net_58215;
  wire net_58216;
  wire net_58221;
  wire net_58223;
  wire net_58233;
  wire net_58236;
  wire net_58241;
  wire net_58243;
  wire net_58250;
  wire net_58251;
  wire net_58253;
  wire net_58254;
  wire net_58264;
  wire net_58268;
  wire net_58270;
  wire net_58273;
  wire net_58274;
  wire net_58275;
  wire net_58284;
  wire net_58285;
  wire net_58296;
  wire net_58298;
  wire net_58307;
  wire net_58308;
  wire net_58313;
  wire net_58314;
  wire net_58319;
  wire net_58320;
  wire net_58321;
  wire net_58322;
  wire net_58325;
  wire net_58327;
  wire net_58329;
  wire net_58330;
  wire net_58331;
  wire net_58332;
  wire net_58333;
  wire net_58334;
  wire net_58335;
  wire net_58336;
  wire net_58338;
  wire net_58339;
  wire net_58346;
  wire net_58350;
  wire net_58354;
  wire net_58355;
  wire net_58357;
  wire net_58358;
  wire net_58361;
  wire net_58363;
  wire net_58365;
  wire net_58367;
  wire net_58373;
  wire net_58375;
  wire net_58378;
  wire net_58380;
  wire net_58385;
  wire net_58386;
  wire net_58387;
  wire net_58388;
  wire net_58393;
  wire net_58396;
  wire net_58407;
  wire net_58412;
  wire net_58413;
  wire net_58415;
  wire net_58419;
  wire net_58427;
  wire net_58431;
  wire net_58436;
  wire net_58444;
  wire net_58449;
  wire net_58453;
  wire net_58454;
  wire net_58456;
  wire net_58457;
  wire net_58458;
  wire net_58459;
  wire net_58460;
  wire net_58461;
  wire net_58462;
  wire net_58467;
  wire net_58481;
  wire net_58483;
  wire net_58486;
  wire net_58488;
  wire net_58489;
  wire net_58496;
  wire net_58499;
  wire net_58500;
  wire net_58501;
  wire net_58503;
  wire net_58504;
  wire net_58506;
  wire net_58507;
  wire net_58509;
  wire net_58510;
  wire net_58511;
  wire net_58514;
  wire net_58516;
  wire net_58522;
  wire net_58527;
  wire net_58531;
  wire net_58534;
  wire net_58536;
  wire net_58537;
  wire net_58540;
  wire net_58542;
  wire net_58543;
  wire net_58544;
  wire net_58546;
  wire net_58548;
  wire net_58549;
  wire net_58550;
  wire net_58552;
  wire net_58554;
  wire net_58555;
  wire net_58556;
  wire net_58558;
  wire net_58560;
  wire net_58561;
  wire net_58562;
  wire net_58564;
  wire net_58566;
  wire net_58567;
  wire net_58568;
  wire net_58570;
  wire net_58572;
  wire net_58573;
  wire net_58574;
  wire net_58576;
  wire net_58577;
  wire net_58578;
  wire net_58579;
  wire net_58580;
  wire net_58582;
  wire net_58592;
  wire net_58596;
  wire net_58600;
  wire net_58603;
  wire net_58604;
  wire net_58605;
  wire net_58610;
  wire net_58614;
  wire net_58620;
  wire net_58621;
  wire net_58626;
  wire net_58630;
  wire net_58633;
  wire net_58646;
  wire net_58651;
  wire net_58653;
  wire net_58654;
  wire net_58655;
  wire net_58661;
  wire net_58665;
  wire net_58672;
  wire net_58685;
  wire net_58690;
  wire net_58697;
  wire net_58699;
  wire net_58700;
  wire net_58705;
  wire net_58713;
  wire net_58716;
  wire net_58717;
  wire net_58720;
  wire net_58742;
  wire net_58743;
  wire net_58745;
  wire net_58747;
  wire net_58748;
  wire net_58750;
  wire net_58751;
  wire net_58752;
  wire net_58753;
  wire net_58754;
  wire net_58756;
  wire net_58761;
  wire net_58764;
  wire net_58765;
  wire net_58768;
  wire net_58769;
  wire net_58770;
  wire net_58775;
  wire net_58776;
  wire net_58777;
  wire net_58781;
  wire net_58782;
  wire net_58783;
  wire net_58787;
  wire net_58788;
  wire net_58789;
  wire net_58790;
  wire net_58794;
  wire net_58795;
  wire net_58796;
  wire net_58806;
  wire net_58807;
  wire net_58808;
  wire net_58811;
  wire net_58812;
  wire net_58813;
  wire net_58814;
  wire net_58817;
  wire net_58818;
  wire net_58819;
  wire net_58820;
  wire net_58821;
  wire net_58822;
  wire net_58823;
  wire net_58847;
  wire net_58883;
  wire net_58884;
  wire net_58889;
  wire net_58892;
  wire net_58896;
  wire net_58916;
  wire net_58917;
  wire net_58918;
  wire net_58919;
  wire net_58944;
  wire net_58945;
  wire net_58946;
  wire net_60411;
  wire net_60431;
  wire net_60530;
  wire net_60590;
  wire net_60627;
  wire net_60676;
  wire net_60683;
  wire net_60684;
  wire net_60688;
  wire net_60689;
  wire net_60701;
  wire net_60705;
  wire net_60729;
  wire net_60731;
  wire net_60774;
  wire net_60784;
  wire net_60807;
  wire net_60808;
  wire net_60810;
  wire net_60811;
  wire net_60812;
  wire net_60813;
  wire net_60814;
  wire net_60815;
  wire net_60816;
  wire net_60833;
  wire net_60834;
  wire net_60835;
  wire net_60837;
  wire net_60842;
  wire net_60844;
  wire net_60850;
  wire net_60852;
  wire net_60860;
  wire net_60866;
  wire net_60870;
  wire net_60874;
  wire net_60876;
  wire net_60878;
  wire net_60880;
  wire net_60886;
  wire net_60890;
  wire net_60892;
  wire net_60895;
  wire net_60901;
  wire net_60904;
  wire net_60908;
  wire net_60909;
  wire net_60914;
  wire net_60915;
  wire net_60921;
  wire net_60922;
  wire net_60926;
  wire net_60930;
  wire net_60931;
  wire net_60932;
  wire net_60933;
  wire net_60934;
  wire net_60935;
  wire net_60936;
  wire net_60937;
  wire net_60938;
  wire net_60939;
  wire net_60952;
  wire net_60956;
  wire net_60958;
  wire net_60959;
  wire net_60960;
  wire net_60961;
  wire net_60964;
  wire net_60965;
  wire net_60966;
  wire net_60967;
  wire net_60973;
  wire net_60978;
  wire net_60982;
  wire net_60983;
  wire net_60988;
  wire net_60991;
  wire net_60993;
  wire net_60998;
  wire net_61001;
  wire net_61006;
  wire net_61007;
  wire net_61013;
  wire net_61015;
  wire net_61018;
  wire net_61020;
  wire net_61025;
  wire net_61027;
  wire net_61032;
  wire net_61033;
  wire net_61036;
  wire net_61039;
  wire net_61042;
  wire net_61044;
  wire net_61049;
  wire net_61051;
  wire net_61053;
  wire net_61054;
  wire net_61056;
  wire net_61057;
  wire net_61058;
  wire net_61059;
  wire net_61060;
  wire net_61061;
  wire net_61062;
  wire net_61079;
  wire net_61081;
  wire net_61085;
  wire net_61096;
  wire net_61097;
  wire net_61098;
  wire net_61099;
  wire net_61100;
  wire net_61102;
  wire net_61104;
  wire net_61106;
  wire net_61107;
  wire net_61108;
  wire net_61109;
  wire net_61111;
  wire net_61112;
  wire net_61114;
  wire net_61115;
  wire net_61116;
  wire net_61117;
  wire net_61118;
  wire net_61121;
  wire net_61122;
  wire net_61123;
  wire net_61124;
  wire net_61125;
  wire net_61127;
  wire net_61129;
  wire net_61130;
  wire net_61131;
  wire net_61132;
  wire net_61135;
  wire net_61136;
  wire net_61137;
  wire net_61138;
  wire net_61147;
  wire net_61148;
  wire net_61149;
  wire net_61150;
  wire net_61153;
  wire net_61154;
  wire net_61155;
  wire net_61156;
  wire net_61159;
  wire net_61160;
  wire net_61161;
  wire net_61162;
  wire net_61165;
  wire net_61166;
  wire net_61167;
  wire net_61168;
  wire net_61171;
  wire net_61172;
  wire net_61173;
  wire net_61174;
  wire net_61175;
  wire net_61176;
  wire net_61177;
  wire net_61178;
  wire net_61179;
  wire net_61180;
  wire net_61181;
  wire net_61182;
  wire net_61183;
  wire net_61184;
  wire net_61185;
  wire net_61194;
  wire net_61201;
  wire net_61204;
  wire net_61205;
  wire net_61208;
  wire net_61212;
  wire net_61213;
  wire net_61234;
  wire net_61241;
  wire net_61242;
  wire net_61246;
  wire net_61266;
  wire net_61272;
  wire net_61276;
  wire net_61290;
  wire net_61299;
  wire net_61300;
  wire net_61301;
  wire net_61302;
  wire net_61305;
  wire net_61316;
  wire net_61320;
  wire net_61322;
  wire net_61324;
  wire net_61325;
  wire net_61335;
  wire net_61336;
  wire net_61345;
  wire net_61347;
  wire net_61355;
  wire net_61366;
  wire net_61382;
  wire net_61390;
  wire net_61395;
  wire net_61400;
  wire net_61422;
  wire net_61423;
  wire net_61425;
  wire net_61426;
  wire net_61428;
  wire net_61429;
  wire net_61430;
  wire net_61431;
  wire net_61432;
  wire net_61438;
  wire net_61439;
  wire net_61443;
  wire net_61452;
  wire net_61459;
  wire net_61468;
  wire net_61469;
  wire net_61475;
  wire net_61476;
  wire net_61485;
  wire net_61492;
  wire net_61496;
  wire net_61498;
  wire net_61506;
  wire net_61513;
  wire net_61519;
  wire net_61524;
  wire net_61536;
  wire net_61544;
  wire net_61545;
  wire net_61547;
  wire net_61548;
  wire net_61549;
  wire net_61550;
  wire net_61551;
  wire net_61552;
  wire net_61553;
  wire net_61554;
  wire net_61571;
  wire net_61572;
  wire net_61573;
  wire net_61574;
  wire net_61576;
  wire net_61577;
  wire net_61578;
  wire net_61588;
  wire net_61594;
  wire net_61596;
  wire net_61597;
  wire net_61602;
  wire net_61606;
  wire net_61607;
  wire net_61610;
  wire net_61614;
  wire net_61622;
  wire net_61626;
  wire net_61627;
  wire net_61628;
  wire net_61630;
  wire net_61632;
  wire net_61633;
  wire net_61634;
  wire net_61636;
  wire net_61639;
  wire net_61641;
  wire net_61642;
  wire net_61657;
  wire net_61664;
  wire net_61666;
  wire net_61667;
  wire net_61668;
  wire net_61669;
  wire net_61671;
  wire net_61672;
  wire net_61673;
  wire net_61674;
  wire net_61675;
  wire net_61676;
  wire net_61677;
  wire net_61682;
  wire net_61686;
  wire net_61702;
  wire net_61713;
  wire net_61714;
  wire net_61720;
  wire net_61723;
  wire net_61724;
  wire net_61725;
  wire net_61731;
  wire net_61733;
  wire net_61734;
  wire net_61736;
  wire net_61737;
  wire net_61742;
  wire net_61744;
  wire net_61746;
  wire net_61747;
  wire net_61751;
  wire net_61752;
  wire net_61753;
  wire net_61756;
  wire net_61765;
  wire net_61769;
  wire net_61776;
  wire net_61780;
  wire net_61788;
  wire net_61791;
  wire net_61792;
  wire net_61795;
  wire net_61796;
  wire net_61799;
  wire net_61800;
  wire net_61805;
  wire net_61812;
  wire net_61823;
  wire net_61825;
  wire net_61826;
  wire net_61841;
  wire net_61843;
  wire net_61849;
  wire net_61851;
  wire net_61852;
  wire net_61854;
  wire net_61857;
  wire net_61864;
  wire net_61865;
  wire net_61869;
  wire net_61870;
  wire net_61874;
  wire net_61882;
  wire net_61887;
  wire net_61891;
  wire net_61899;
  wire net_61903;
  wire net_61910;
  wire net_61914;
  wire net_61915;
  wire net_61917;
  wire net_61918;
  wire net_61919;
  wire net_61920;
  wire net_61921;
  wire net_61922;
  wire net_61923;
  wire net_61929;
  wire net_61939;
  wire net_61948;
  wire net_61951;
  wire net_61962;
  wire net_61968;
  wire net_61975;
  wire net_61976;
  wire net_61982;
  wire net_61985;
  wire net_61986;
  wire net_61987;
  wire net_61989;
  wire net_61991;
  wire net_61992;
  wire net_61995;
  wire net_61997;
  wire net_61999;
  wire net_62001;
  wire net_62004;
  wire net_62005;
  wire net_62007;
  wire net_62010;
  wire net_62011;
  wire net_62013;
  wire net_62015;
  wire net_62017;
  wire net_62019;
  wire net_62021;
  wire net_62023;
  wire net_62025;
  wire net_62027;
  wire net_62029;
  wire net_62035;
  wire net_62037;
  wire net_62038;
  wire net_62040;
  wire net_62041;
  wire net_62042;
  wire net_62043;
  wire net_62044;
  wire net_62045;
  wire net_62046;
  wire net_62052;
  wire net_62058;
  wire net_62062;
  wire net_62066;
  wire net_62068;
  wire net_62073;
  wire net_62081;
  wire net_62082;
  wire net_62083;
  wire net_62085;
  wire net_62090;
  wire net_62091;
  wire net_62092;
  wire net_62093;
  wire net_62096;
  wire net_62097;
  wire net_62107;
  wire net_62109;
  wire net_62115;
  wire net_62119;
  wire net_62121;
  wire net_62127;
  wire net_62128;
  wire net_62131;
  wire net_62133;
  wire net_62138;
  wire net_62140;
  wire net_62144;
  wire net_62145;
  wire net_62150;
  wire net_62152;
  wire net_62156;
  wire net_62158;
  wire net_62159;
  wire net_62160;
  wire net_62161;
  wire net_62162;
  wire net_62163;
  wire net_62164;
  wire net_62165;
  wire net_62166;
  wire net_62167;
  wire net_62168;
  wire net_62169;
  wire net_62174;
  wire net_62175;
  wire net_62179;
  wire net_62180;
  wire net_62181;
  wire net_62187;
  wire net_62193;
  wire net_62197;
  wire net_62212;
  wire net_62213;
  wire net_62214;
  wire net_62228;
  wire net_62232;
  wire net_62233;
  wire net_62236;
  wire net_62245;
  wire net_62250;
  wire net_62256;
  wire net_62261;
  wire net_62272;
  wire net_62280;
  wire net_62283;
  wire net_62284;
  wire net_62285;
  wire net_62286;
  wire net_62287;
  wire net_62288;
  wire net_62289;
  wire net_62290;
  wire net_62291;
  wire net_62292;
  wire net_62298;
  wire net_62326;
  wire net_62327;
  wire net_62331;
  wire net_62333;
  wire net_62335;
  wire net_62337;
  wire net_62342;
  wire net_62345;
  wire net_62347;
  wire net_62348;
  wire net_62351;
  wire net_62352;
  wire net_62353;
  wire net_62355;
  wire net_62356;
  wire net_62361;
  wire net_62364;
  wire net_62366;
  wire net_62367;
  wire net_62368;
  wire net_62370;
  wire net_62372;
  wire net_62373;
  wire net_62374;
  wire net_62376;
  wire net_62378;
  wire net_62379;
  wire net_62380;
  wire net_62382;
  wire net_62384;
  wire net_62385;
  wire net_62386;
  wire net_62388;
  wire net_62390;
  wire net_62391;
  wire net_62392;
  wire net_62394;
  wire net_62396;
  wire net_62397;
  wire net_62398;
  wire net_62400;
  wire net_62402;
  wire net_62403;
  wire net_62404;
  wire net_62406;
  wire net_62407;
  wire net_62408;
  wire net_62409;
  wire net_62410;
  wire net_62411;
  wire net_62412;
  wire net_62413;
  wire net_62414;
  wire net_62415;
  wire net_62444;
  wire net_62449;
  wire net_62466;
  wire net_62467;
  wire net_62468;
  wire net_62470;
  wire net_62480;
  wire net_62481;
  wire net_62483;
  wire net_62484;
  wire net_62485;
  wire net_62491;
  wire net_62496;
  wire net_62506;
  wire net_62507;
  wire net_62509;
  wire net_62529;
  wire net_62530;
  wire net_62531;
  wire net_62543;
  wire net_62547;
  wire net_62548;
  wire net_62555;
  wire net_62575;
  wire net_62582;
  wire net_62583;
  wire net_62592;
  wire net_62597;
  wire net_62629;
  wire net_62630;
  wire net_62631;
  wire net_62632;
  wire net_62651;
  wire net_62652;
  wire net_62653;
  wire net_64205;
  wire net_64225;
  wire net_64260;
  wire net_64262;
  wire net_64354;
  wire net_64358;
  wire net_64365;
  wire net_64408;
  wire net_64424;
  wire net_64440;
  wire net_64488;
  wire net_64514;
  wire net_64515;
  wire net_64517;
  wire net_64518;
  wire net_64519;
  wire net_64520;
  wire net_64521;
  wire net_64529;
  wire net_64534;
  wire net_64560;
  wire net_64564;
  wire net_64568;
  wire net_64569;
  wire net_64580;
  wire net_64585;
  wire net_64586;
  wire net_64603;
  wire net_64604;
  wire net_64605;
  wire net_64606;
  wire net_64610;
  wire net_64612;
  wire net_64637;
  wire net_64638;
  wire net_64639;
  wire net_64640;
  wire net_64641;
  wire net_64642;
  wire net_64643;
  wire net_64644;
  wire net_64645;
  wire net_64646;
  wire net_64647;
  wire net_64658;
  wire net_64660;
  wire net_64665;
  wire net_64666;
  wire net_64674;
  wire net_64685;
  wire net_64688;
  wire net_64692;
  wire net_64693;
  wire net_64695;
  wire net_64696;
  wire net_64697;
  wire net_64698;
  wire net_64699;
  wire net_64700;
  wire net_64701;
  wire net_64702;
  wire net_64703;
  wire net_64705;
  wire net_64711;
  wire net_64712;
  wire net_64713;
  wire net_64715;
  wire net_64716;
  wire net_64719;
  wire net_64721;
  wire net_64722;
  wire net_64723;
  wire net_64725;
  wire net_64727;
  wire net_64728;
  wire net_64729;
  wire net_64731;
  wire net_64733;
  wire net_64734;
  wire net_64735;
  wire net_64737;
  wire net_64739;
  wire net_64740;
  wire net_64741;
  wire net_64743;
  wire net_64745;
  wire net_64746;
  wire net_64747;
  wire net_64749;
  wire net_64751;
  wire net_64752;
  wire net_64753;
  wire net_64755;
  wire net_64757;
  wire net_64758;
  wire net_64759;
  wire net_64763;
  wire net_64764;
  wire net_64765;
  wire net_64766;
  wire net_64768;
  wire net_64769;
  wire net_64770;
  wire net_64771;
  wire net_64792;
  wire net_64796;
  wire net_64798;
  wire net_64799;
  wire net_64805;
  wire net_64812;
  wire net_64817;
  wire net_64820;
  wire net_64822;
  wire net_64823;
  wire net_64826;
  wire net_64829;
  wire net_64830;
  wire net_64834;
  wire net_64835;
  wire net_64836;
  wire net_64838;
  wire net_64839;
  wire net_64840;
  wire net_64842;
  wire net_64844;
  wire net_64845;
  wire net_64846;
  wire net_64848;
  wire net_64850;
  wire net_64851;
  wire net_64852;
  wire net_64858;
  wire net_64861;
  wire net_64868;
  wire net_64870;
  wire net_64876;
  wire net_64881;
  wire net_64884;
  wire net_64885;
  wire net_64888;
  wire net_64890;
  wire net_64891;
  wire net_64892;
  wire net_64893;
  wire net_64911;
  wire net_64912;
  wire net_64913;
  wire net_64920;
  wire net_64929;
  wire net_64931;
  wire net_64932;
  wire net_64933;
  wire net_64938;
  wire net_64941;
  wire net_64946;
  wire net_64952;
  wire net_64956;
  wire net_64959;
  wire net_64961;
  wire net_64962;
  wire net_64965;
  wire net_64968;
  wire net_64969;
  wire net_64971;
  wire net_64974;
  wire net_64975;
  wire net_64977;
  wire net_64979;
  wire net_64981;
  wire net_64983;
  wire net_64986;
  wire net_64987;
  wire net_64989;
  wire net_64991;
  wire net_64993;
  wire net_64995;
  wire net_64998;
  wire net_64999;
  wire net_65001;
  wire net_65004;
  wire net_65005;
  wire net_65007;
  wire net_65008;
  wire net_65016;
  wire net_65020;
  wire net_65026;
  wire net_65037;
  wire net_65042;
  wire net_65045;
  wire net_65050;
  wire net_65052;
  wire net_65053;
  wire net_65054;
  wire net_65062;
  wire net_65065;
  wire net_65070;
  wire net_65073;
  wire net_65082;
  wire net_65085;
  wire net_65086;
  wire net_65088;
  wire net_65090;
  wire net_65092;
  wire net_65094;
  wire net_65096;
  wire net_65098;
  wire net_65100;
  wire net_65103;
  wire net_65104;
  wire net_65110;
  wire net_65116;
  wire net_65121;
  wire net_65122;
  wire net_65126;
  wire net_65130;
  wire net_65131;
  wire net_65133;
  wire net_65134;
  wire net_65138;
  wire net_65144;
  wire net_65148;
  wire net_65150;
  wire net_65165;
  wire net_65167;
  wire net_65176;
  wire net_65180;
  wire net_65185;
  wire net_65186;
  wire net_65207;
  wire net_65212;
  wire net_65214;
  wire net_65232;
  wire net_65253;
  wire net_65254;
  wire net_65259;
  wire net_65262;
  wire net_65265;
  wire net_65277;
  wire net_65279;
  wire net_65284;
  wire net_65288;
  wire net_65290;
  wire net_65303;
  wire net_65304;
  wire net_65307;
  wire net_65310;
  wire net_65319;
  wire net_65327;
  wire net_65337;
  wire net_65344;
  wire net_65356;
  wire net_65362;
  wire net_65366;
  wire net_65372;
  wire net_65376;
  wire net_65377;
  wire net_65378;
  wire net_65379;
  wire net_65380;
  wire net_65381;
  wire net_65382;
  wire net_65383;
  wire net_65385;
  wire net_65392;
  wire net_65402;
  wire net_65405;
  wire net_65406;
  wire net_65408;
  wire net_65410;
  wire net_65411;
  wire net_65421;
  wire net_65423;
  wire net_65427;
  wire net_65428;
  wire net_65436;
  wire net_65438;
  wire net_65439;
  wire net_65444;
  wire net_65445;
  wire net_65446;
  wire net_65454;
  wire net_65455;
  wire net_65458;
  wire net_65461;
  wire net_65464;
  wire net_65465;
  wire net_65470;
  wire net_65472;
  wire net_65477;
  wire net_65478;
  wire net_65482;
  wire net_65485;
  wire net_65489;
  wire net_65491;
  wire net_65494;
  wire net_65495;
  wire net_65499;
  wire net_65500;
  wire net_65502;
  wire net_65503;
  wire net_65504;
  wire net_65505;
  wire net_65506;
  wire net_65507;
  wire net_65508;
  wire net_65511;
  wire net_65517;
  wire net_65521;
  wire net_65528;
  wire net_65530;
  wire net_65532;
  wire net_65543;
  wire net_65544;
  wire net_65546;
  wire net_65547;
  wire net_65555;
  wire net_65562;
  wire net_65565;
  wire net_65567;
  wire net_65568;
  wire net_65569;
  wire net_65571;
  wire net_65572;
  wire net_65573;
  wire net_65574;
  wire net_65576;
  wire net_65577;
  wire net_65580;
  wire net_65581;
  wire net_65582;
  wire net_65583;
  wire net_65584;
  wire net_65586;
  wire net_65587;
  wire net_65588;
  wire net_65589;
  wire net_65590;
  wire net_65592;
  wire net_65593;
  wire net_65594;
  wire net_65595;
  wire net_65596;
  wire net_65598;
  wire net_65599;
  wire net_65600;
  wire net_65601;
  wire net_65602;
  wire net_65608;
  wire net_65611;
  wire net_65612;
  wire net_65613;
  wire net_65618;
  wire net_65620;
  wire net_65621;
  wire net_65622;
  wire net_65623;
  wire net_65624;
  wire net_65625;
  wire net_65626;
  wire net_65627;
  wire net_65628;
  wire net_65629;
  wire net_65630;
  wire net_65631;
  wire net_65636;
  wire net_65646;
  wire net_65651;
  wire net_65667;
  wire net_65668;
  wire net_65670;
  wire net_65672;
  wire net_65673;
  wire net_65674;
  wire net_65677;
  wire net_65678;
  wire net_65679;
  wire net_65680;
  wire net_65682;
  wire net_65686;
  wire net_65690;
  wire net_65694;
  wire net_65710;
  wire net_65711;
  wire net_65712;
  wire net_65713;
  wire net_65716;
  wire net_65717;
  wire net_65718;
  wire net_65719;
  wire net_65734;
  wire net_65735;
  wire net_65736;
  wire net_65737;
  wire net_65740;
  wire net_65741;
  wire net_65742;
  wire net_65743;
  wire net_65744;
  wire net_65745;
  wire net_65748;
  wire net_65749;
  wire net_65750;
  wire net_65751;
  wire net_65752;
  wire net_65753;
  wire net_65777;
  wire net_65781;
  wire net_65790;
  wire net_65792;
  wire net_65796;
  wire net_65797;
  wire net_65799;
  wire net_65800;
  wire net_65806;
  wire net_65807;
  wire net_65810;
  wire net_65812;
  wire net_65813;
  wire net_65814;
  wire net_65815;
  wire net_65816;
  wire net_65819;
  wire net_65820;
  wire net_65822;
  wire net_65823;
  wire net_65826;
  wire net_65828;
  wire net_65829;
  wire net_65830;
  wire net_65832;
  wire net_65834;
  wire net_65835;
  wire net_65836;
  wire net_65838;
  wire net_65840;
  wire net_65841;
  wire net_65842;
  wire net_65844;
  wire net_65846;
  wire net_65847;
  wire net_65848;
  wire net_65850;
  wire net_65852;
  wire net_65853;
  wire net_65854;
  wire net_65860;
  wire net_65864;
  wire net_65866;
  wire net_65867;
  wire net_65868;
  wire net_65869;
  wire net_65870;
  wire net_65871;
  wire net_65872;
  wire net_65873;
  wire net_65874;
  wire net_65875;
  wire net_65876;
  wire net_65877;
  wire net_65884;
  wire net_65894;
  wire net_65899;
  wire net_65901;
  wire net_65903;
  wire net_65904;
  wire net_65905;
  wire net_65911;
  wire net_65912;
  wire net_65913;
  wire net_65917;
  wire net_65919;
  wire net_65923;
  wire net_65924;
  wire net_65925;
  wire net_65926;
  wire net_65930;
  wire net_65933;
  wire net_65934;
  wire net_65935;
  wire net_65937;
  wire net_65938;
  wire net_65940;
  wire net_65943;
  wire net_65945;
  wire net_65946;
  wire net_65949;
  wire net_65951;
  wire net_65952;
  wire net_65953;
  wire net_65955;
  wire net_65957;
  wire net_65958;
  wire net_65959;
  wire net_65961;
  wire net_65963;
  wire net_65964;
  wire net_65965;
  wire net_65967;
  wire net_65969;
  wire net_65970;
  wire net_65971;
  wire net_65973;
  wire net_65975;
  wire net_65976;
  wire net_65977;
  wire net_65979;
  wire net_65981;
  wire net_65982;
  wire net_65983;
  wire net_65985;
  wire net_65987;
  wire net_65988;
  wire net_65989;
  wire net_65993;
  wire net_65994;
  wire net_65995;
  wire net_65996;
  wire net_65997;
  wire net_65998;
  wire net_65999;
  wire net_66000;
  wire net_66013;
  wire net_66015;
  wire net_66017;
  wire net_66019;
  wire net_66021;
  wire net_66025;
  wire net_66029;
  wire net_66040;
  wire net_66041;
  wire net_66049;
  wire net_66050;
  wire net_66051;
  wire net_66054;
  wire net_66063;
  wire net_66064;
  wire net_66067;
  wire net_66069;
  wire net_66070;
  wire net_66075;
  wire net_66080;
  wire net_66086;
  wire net_66092;
  wire net_66100;
  wire net_66105;
  wire net_66112;
  wire net_66114;
  wire net_66115;
  wire net_66117;
  wire net_66118;
  wire net_66119;
  wire net_66120;
  wire net_66121;
  wire net_66122;
  wire net_66130;
  wire net_66141;
  wire net_66142;
  wire net_66160;
  wire net_66161;
  wire net_66162;
  wire net_66164;
  wire net_66165;
  wire net_66167;
  wire net_66169;
  wire net_66171;
  wire net_66172;
  wire net_66176;
  wire net_66180;
  wire net_66185;
  wire net_66187;
  wire net_66188;
  wire net_66190;
  wire net_66191;
  wire net_66192;
  wire net_66193;
  wire net_66196;
  wire net_66197;
  wire net_66198;
  wire net_66199;
  wire net_66202;
  wire net_66203;
  wire net_66204;
  wire net_66205;
  wire net_66209;
  wire net_66210;
  wire net_66215;
  wire net_66216;
  wire net_66221;
  wire net_66223;
  wire net_66226;
  wire net_66227;
  wire net_66228;
  wire net_66229;
  wire net_66234;
  wire net_66235;
  wire net_66236;
  wire net_66237;
  wire net_66238;
  wire net_66239;
  wire net_66240;
  wire net_66242;
  wire net_66243;
  wire net_66244;
  wire net_66245;
  wire net_66246;
  wire net_66253;
  wire net_66261;
  wire net_66280;
  wire net_66282;
  wire net_66283;
  wire net_66284;
  wire net_66293;
  wire net_66297;
  wire net_66299;
  wire net_66302;
  wire net_66303;
  wire net_66304;
  wire net_66305;
  wire net_66308;
  wire net_66310;
  wire net_66314;
  wire net_66315;
  wire net_66319;
  wire net_66321;
  wire net_66325;
  wire net_66326;
  wire net_66327;
  wire net_66328;
  wire net_66331;
  wire net_66332;
  wire net_66338;
  wire net_66340;
  wire net_66343;
  wire net_66345;
  wire net_66349;
  wire net_66350;
  wire net_66355;
  wire net_66356;
  wire net_66357;
  wire net_66358;
  wire net_66359;
  wire net_66360;
  wire net_66361;
  wire net_66368;
  wire net_66379;
  wire net_66391;
  wire net_66393;
  wire net_66414;
  wire net_66425;
  wire net_66438;
  wire net_66482;
  wire net_66483;
  wire net_66484;
  wire net_68006;
  wire net_68009;
  wire net_68021;
  wire net_68025;
  wire net_68185;
  wire net_68193;
  wire net_68248;
  wire net_68281;
  wire net_68292;
  wire net_68299;
  wire net_68341;
  wire net_68345;
  wire net_68346;
  wire net_68348;
  wire net_68349;
  wire net_68350;
  wire net_68351;
  wire net_68352;
  wire net_68353;
  wire net_68354;
  wire net_68355;
  wire net_68360;
  wire net_68361;
  wire net_68363;
  wire net_68391;
  wire net_68392;
  wire net_68400;
  wire net_68409;
  wire net_68413;
  wire net_68424;
  wire net_68430;
  wire net_68436;
  wire net_68440;
  wire net_68446;
  wire net_68469;
  wire net_68470;
  wire net_68472;
  wire net_68473;
  wire net_68474;
  wire net_68475;
  wire net_68476;
  wire net_68477;
  wire net_68478;
  wire net_68486;
  wire net_68488;
  wire net_68492;
  wire net_68496;
  wire net_68503;
  wire net_68504;
  wire net_68515;
  wire net_68520;
  wire net_68522;
  wire net_68523;
  wire net_68525;
  wire net_68526;
  wire net_68527;
  wire net_68535;
  wire net_68546;
  wire net_68553;
  wire net_68560;
  wire net_68566;
  wire net_68572;
  wire net_68578;
  wire net_68583;
  wire net_68589;
  wire net_68592;
  wire net_68593;
  wire net_68594;
  wire net_68595;
  wire net_68596;
  wire net_68597;
  wire net_68598;
  wire net_68599;
  wire net_68600;
  wire net_68601;
  wire net_68618;
  wire net_68620;
  wire net_68622;
  wire net_68624;
  wire net_68638;
  wire net_68642;
  wire net_68643;
  wire net_68644;
  wire net_68646;
  wire net_68653;
  wire net_68666;
  wire net_68670;
  wire net_68674;
  wire net_68682;
  wire net_68687;
  wire net_68698;
  wire net_68706;
  wire net_68712;
  wire net_68715;
  wire net_68716;
  wire net_68717;
  wire net_68718;
  wire net_68720;
  wire net_68721;
  wire net_68722;
  wire net_68723;
  wire net_68724;
  wire net_68730;
  wire net_68732;
  wire net_68734;
  wire net_68736;
  wire net_68738;
  wire net_68743;
  wire net_68752;
  wire net_68764;
  wire net_68771;
  wire net_68779;
  wire net_68783;
  wire net_68785;
  wire net_68805;
  wire net_68815;
  wire net_68822;
  wire net_68827;
  wire net_68835;
  wire net_68838;
  wire net_68839;
  wire net_68841;
  wire net_68842;
  wire net_68843;
  wire net_68844;
  wire net_68845;
  wire net_68846;
  wire net_68847;
  wire net_68850;
  wire net_68859;
  wire net_68865;
  wire net_68869;
  wire net_68875;
  wire net_68888;
  wire net_68899;
  wire net_68958;
  wire net_68960;
  wire net_68961;
  wire net_68962;
  wire net_68963;
  wire net_68964;
  wire net_68967;
  wire net_68968;
  wire net_68970;
  wire net_68980;
  wire net_68984;
  wire net_68986;
  wire net_68987;
  wire net_68989;
  wire net_68993;
  wire net_68995;
  wire net_68996;
  wire net_68997;
  wire net_69005;
  wire net_69006;
  wire net_69009;
  wire net_69013;
  wire net_69014;
  wire net_69019;
  wire net_69020;
  wire net_69022;
  wire net_69024;
  wire net_69028;
  wire net_69030;
  wire net_69032;
  wire net_69043;
  wire net_69044;
  wire net_69045;
  wire net_69046;
  wire net_69049;
  wire net_69050;
  wire net_69051;
  wire net_69052;
  wire net_69073;
  wire net_69074;
  wire net_69075;
  wire net_69076;
  wire net_69083;
  wire net_69084;
  wire net_69086;
  wire net_69087;
  wire net_69089;
  wire net_69091;
  wire net_69092;
  wire net_69107;
  wire net_69128;
  wire net_69131;
  wire net_69185;
  wire net_69203;
  wire net_69207;
  wire net_69208;
  wire net_69210;
  wire net_69211;
  wire net_69212;
  wire net_69213;
  wire net_69214;
  wire net_69215;
  wire net_69216;
  wire net_69230;
  wire net_69254;
  wire net_69258;
  wire net_69263;
  wire net_69265;
  wire net_69269;
  wire net_69270;
  wire net_69280;
  wire net_69286;
  wire net_69292;
  wire net_69295;
  wire net_69303;
  wire net_69308;
  wire net_69316;
  wire net_69326;
  wire net_69330;
  wire net_69331;
  wire net_69332;
  wire net_69333;
  wire net_69334;
  wire net_69335;
  wire net_69336;
  wire net_69337;
  wire net_69338;
  wire net_69339;
  wire net_69357;
  wire net_69358;
  wire net_69367;
  wire net_69373;
  wire net_69374;
  wire net_69378;
  wire net_69380;
  wire net_69381;
  wire net_69384;
  wire net_69385;
  wire net_69386;
  wire net_69388;
  wire net_69389;
  wire net_69391;
  wire net_69395;
  wire net_69397;
  wire net_69399;
  wire net_69402;
  wire net_69403;
  wire net_69405;
  wire net_69407;
  wire net_69408;
  wire net_69411;
  wire net_69413;
  wire net_69414;
  wire net_69415;
  wire net_69417;
  wire net_69419;
  wire net_69420;
  wire net_69421;
  wire net_69423;
  wire net_69425;
  wire net_69426;
  wire net_69427;
  wire net_69429;
  wire net_69431;
  wire net_69433;
  wire net_69436;
  wire net_69437;
  wire net_69438;
  wire net_69439;
  wire net_69442;
  wire net_69445;
  wire net_69448;
  wire net_69449;
  wire net_69452;
  wire net_69453;
  wire net_69454;
  wire net_69455;
  wire net_69456;
  wire net_69457;
  wire net_69458;
  wire net_69459;
  wire net_69461;
  wire net_69462;
  wire net_69499;
  wire net_69509;
  wire net_69515;
  wire net_69518;
  wire net_69521;
  wire net_69522;
  wire net_69525;
  wire net_69526;
  wire net_69532;
  wire net_69535;
  wire net_69541;
  wire net_69549;
  wire net_69555;
  wire net_69560;
  wire net_69568;
  wire net_69574;
  wire net_69576;
  wire net_69577;
  wire net_69578;
  wire net_69579;
  wire net_69580;
  wire net_69582;
  wire net_69583;
  wire net_69584;
  wire net_69602;
  wire net_69604;
  wire net_69610;
  wire net_69623;
  wire net_69637;
  wire net_69638;
  wire net_69639;
  wire net_69641;
  wire net_69644;
  wire net_69646;
  wire net_69648;
  wire net_69650;
  wire net_69651;
  wire net_69653;
  wire net_69654;
  wire net_69657;
  wire net_69659;
  wire net_69660;
  wire net_69661;
  wire net_69663;
  wire net_69665;
  wire net_69666;
  wire net_69667;
  wire net_69669;
  wire net_69671;
  wire net_69672;
  wire net_69673;
  wire net_69675;
  wire net_69677;
  wire net_69678;
  wire net_69679;
  wire net_69681;
  wire net_69683;
  wire net_69684;
  wire net_69685;
  wire net_69689;
  wire net_69690;
  wire net_69691;
  wire net_69693;
  wire net_69695;
  wire net_69696;
  wire net_69701;
  wire net_69702;
  wire net_69703;
  wire net_69704;
  wire net_69705;
  wire net_69706;
  wire net_69707;
  wire net_69708;
  wire net_69717;
  wire net_69728;
  wire net_69730;
  wire net_69736;
  wire net_69737;
  wire net_69744;
  wire net_69746;
  wire net_69747;
  wire net_69748;
  wire net_69753;
  wire net_69754;
  wire net_69755;
  wire net_69756;
  wire net_69757;
  wire net_69758;
  wire net_69760;
  wire net_69762;
  wire net_69763;
  wire net_69764;
  wire net_69765;
  wire net_69766;
  wire net_69768;
  wire net_69770;
  wire net_69772;
  wire net_69773;
  wire net_69775;
  wire net_69777;
  wire net_69778;
  wire net_69781;
  wire net_69782;
  wire net_69783;
  wire net_69784;
  wire net_69787;
  wire net_69788;
  wire net_69789;
  wire net_69790;
  wire net_69793;
  wire net_69794;
  wire net_69795;
  wire net_69796;
  wire net_69799;
  wire net_69800;
  wire net_69801;
  wire net_69808;
  wire net_69811;
  wire net_69812;
  wire net_69813;
  wire net_69814;
  wire net_69817;
  wire net_69818;
  wire net_69819;
  wire net_69820;
  wire net_69821;
  wire net_69822;
  wire net_69823;
  wire net_69825;
  wire net_69826;
  wire net_69827;
  wire net_69828;
  wire net_69829;
  wire net_69830;
  wire net_69831;
  wire net_69836;
  wire net_69841;
  wire net_69850;
  wire net_69868;
  wire net_69882;
  wire net_69883;
  wire net_69884;
  wire net_69886;
  wire net_69891;
  wire net_69892;
  wire net_69894;
  wire net_69900;
  wire net_69905;
  wire net_69911;
  wire net_69918;
  wire net_69925;
  wire net_69930;
  wire net_69934;
  wire net_69940;
  wire net_69945;
  wire net_69946;
  wire net_69947;
  wire net_69948;
  wire net_69949;
  wire net_69951;
  wire net_69952;
  wire net_69954;
  wire net_69965;
  wire net_69972;
  wire net_69978;
  wire net_69990;
  wire net_69991;
  wire net_69997;
  wire net_70000;
  wire net_70001;
  wire net_70002;
  wire net_70003;
  wire net_70008;
  wire net_70016;
  wire net_70020;
  wire net_70022;
  wire net_70023;
  wire net_70026;
  wire net_70028;
  wire net_70030;
  wire net_70032;
  wire net_70035;
  wire net_70036;
  wire net_70038;
  wire net_70041;
  wire net_70042;
  wire net_70044;
  wire net_70046;
  wire net_70048;
  wire net_70050;
  wire net_70052;
  wire net_70054;
  wire net_70058;
  wire net_70060;
  wire net_70062;
  wire net_70064;
  wire net_70074;
  wire net_70106;
  wire net_70111;
  wire net_70114;
  wire net_70115;
  wire net_70116;
  wire net_70117;
  wire net_70118;
  wire net_70119;
  wire net_70120;
  wire net_70124;
  wire net_70131;
  wire net_70134;
  wire net_70138;
  wire net_70147;
  wire net_70150;
  wire net_70151;
  wire net_70152;
  wire net_70153;
  wire net_70163;
  wire net_70165;
  wire net_70168;
  wire net_70169;
  wire net_70170;
  wire net_70171;
  wire net_70174;
  wire net_70177;
  wire net_70180;
  wire net_70181;
  wire net_70182;
  wire net_70183;
  wire net_70186;
  wire net_70187;
  wire net_70188;
  wire net_70189;
  wire net_70190;
  wire net_70191;
  wire net_70192;
  wire net_70238;
  wire net_70303;
  wire net_70314;
  wire net_70315;
  wire net_71837;
  wire net_71855;
  wire net_71870;
  wire net_71884;
  wire net_72016;
  wire net_72018;
  wire net_72048;
  wire net_72103;
  wire net_72109;
  wire net_72116;
  wire net_72154;
  wire net_72155;
  wire net_72157;
  wire net_72177;
  wire net_72178;
  wire net_72222;
  wire net_72223;
  wire net_72224;
  wire net_72228;
  wire net_72229;
  wire net_72233;
  wire net_72235;
  wire net_72249;
  wire net_72253;
  wire net_72261;
  wire net_72267;
  wire net_72272;
  wire net_72279;
  wire net_72285;
  wire net_72289;
  wire net_72298;
  wire net_72300;
  wire net_72301;
  wire net_72315;
  wire net_72317;
  wire net_72320;
  wire net_72344;
  wire net_72345;
  wire net_72346;
  wire net_72347;
  wire net_72349;
  wire net_72350;
  wire net_72351;
  wire net_72352;
  wire net_72353;
  wire net_72354;
  wire net_72355;
  wire net_72356;
  wire net_72358;
  wire net_72359;
  wire net_72360;
  wire net_72364;
  wire net_72375;
  wire net_72377;
  wire net_72378;
  wire net_72381;
  wire net_72383;
  wire net_72384;
  wire net_72385;
  wire net_72387;
  wire net_72389;
  wire net_72390;
  wire net_72391;
  wire net_72393;
  wire net_72395;
  wire net_72396;
  wire net_72397;
  wire net_72399;
  wire net_72401;
  wire net_72402;
  wire net_72403;
  wire net_72405;
  wire net_72407;
  wire net_72408;
  wire net_72409;
  wire net_72411;
  wire net_72413;
  wire net_72414;
  wire net_72415;
  wire net_72417;
  wire net_72419;
  wire net_72420;
  wire net_72421;
  wire net_72435;
  wire net_72438;
  wire net_72440;
  wire net_72441;
  wire net_72446;
  wire net_72452;
  wire net_72458;
  wire net_72460;
  wire net_72461;
  wire net_72469;
  wire net_72470;
  wire net_72472;
  wire net_72474;
  wire net_72475;
  wire net_72477;
  wire net_72478;
  wire net_72479;
  wire net_72482;
  wire net_72495;
  wire net_72498;
  wire net_72500;
  wire net_72501;
  wire net_72502;
  wire net_72505;
  wire net_72506;
  wire net_72508;
  wire net_72511;
  wire net_72520;
  wire net_72524;
  wire net_72532;
  wire net_72537;
  wire net_72542;
  wire net_72546;
  wire net_72547;
  wire net_72560;
  wire net_72561;
  wire net_72564;
  wire net_72566;
  wire net_72567;
  wire net_72571;
  wire net_72590;
  wire net_72594;
  wire net_72597;
  wire net_72598;
  wire net_72599;
  wire net_72604;
  wire net_72612;
  wire net_72618;
  wire net_72624;
  wire net_72630;
  wire net_72642;
  wire net_72647;
  wire net_72652;
  wire net_72658;
  wire net_72664;
  wire net_72667;
  wire net_72669;
  wire net_72670;
  wire net_72690;
  wire net_72692;
  wire net_72693;
  wire net_72702;
  wire net_72717;
  wire net_72718;
  wire net_72719;
  wire net_72721;
  wire net_72723;
  wire net_72725;
  wire net_72727;
  wire net_72728;
  wire net_72730;
  wire net_72734;
  wire net_72742;
  wire net_72744;
  wire net_72746;
  wire net_72747;
  wire net_72750;
  wire net_72752;
  wire net_72753;
  wire net_72754;
  wire net_72756;
  wire net_72758;
  wire net_72759;
  wire net_72760;
  wire net_72762;
  wire net_72764;
  wire net_72765;
  wire net_72766;
  wire net_72768;
  wire net_72770;
  wire net_72771;
  wire net_72772;
  wire net_72774;
  wire net_72776;
  wire net_72777;
  wire net_72778;
  wire net_72780;
  wire net_72782;
  wire net_72783;
  wire net_72784;
  wire net_72786;
  wire net_72788;
  wire net_72789;
  wire net_72790;
  wire net_72792;
  wire net_72793;
  wire net_72809;
  wire net_72810;
  wire net_72811;
  wire net_72829;
  wire net_72830;
  wire net_72836;
  wire net_72840;
  wire net_72846;
  wire net_72848;
  wire net_72850;
  wire net_72854;
  wire net_72867;
  wire net_72869;
  wire net_72870;
  wire net_72871;
  wire net_72874;
  wire net_72875;
  wire net_72877;
  wire net_72893;
  wire net_72898;
  wire net_72913;
  wire net_72915;
  wire net_72916;
  wire net_72929;
  wire net_72933;
  wire net_72936;
  wire net_72940;
  wire net_72950;
  wire net_72970;
  wire net_72971;
  wire net_72973;
  wire net_72974;
  wire net_72976;
  wire net_72987;
  wire net_72991;
  wire net_72993;
  wire net_72997;
  wire net_73012;
  wire net_73022;
  wire net_73029;
  wire net_73038;
  wire net_73039;
  wire net_73081;
  wire net_73082;
  wire net_73086;
  wire net_73087;
  wire net_73091;
  wire net_73094;
  wire net_73095;
  wire net_73096;
  wire net_73097;
  wire net_73103;
  wire net_73104;
  wire net_73106;
  wire net_73107;
  wire net_73113;
  wire net_73115;
  wire net_73116;
  wire net_73119;
  wire net_73121;
  wire net_73122;
  wire net_73123;
  wire net_73125;
  wire net_73127;
  wire net_73128;
  wire net_73129;
  wire net_73131;
  wire net_73133;
  wire net_73134;
  wire net_73135;
  wire net_73137;
  wire net_73139;
  wire net_73140;
  wire net_73141;
  wire net_73143;
  wire net_73145;
  wire net_73146;
  wire net_73147;
  wire net_73153;
  wire net_73157;
  wire net_73161;
  wire net_73162;
  wire net_73175;
  wire net_73179;
  wire net_73182;
  wire net_73205;
  wire net_73210;
  wire net_73211;
  wire net_73218;
  wire net_73220;
  wire net_73223;
  wire net_73225;
  wire net_73228;
  wire net_73240;
  wire net_73243;
  wire net_73250;
  wire net_73258;
  wire net_73264;
  wire net_73267;
  wire net_73275;
  wire net_73279;
  wire net_73284;
  wire net_73285;
  wire net_73306;
  wire net_73308;
  wire net_73320;
  wire net_73330;
  wire net_73331;
  wire net_73335;
  wire net_73336;
  wire net_73342;
  wire net_73352;
  wire net_73353;
  wire net_73360;
  wire net_73367;
  wire net_73375;
  wire net_73381;
  wire net_73386;
  wire net_73399;
  wire net_73404;
  wire net_73407;
  wire net_73408;
  wire net_73451;
  wire net_73459;
  wire net_73467;
  wire net_73475;
  wire net_73477;
  wire net_73481;
  wire net_73486;
  wire net_73492;
  wire net_73497;
  wire net_73507;
  wire net_73513;
  wire net_73521;
  wire net_73530;
  wire net_73531;
  wire net_73573;
  wire net_73575;
  wire net_73576;
  wire net_73582;
  wire net_73584;
  wire net_73587;
  wire net_73590;
  wire net_73599;
  wire net_73608;
  wire net_73612;
  wire net_73618;
  wire net_73626;
  wire net_73631;
  wire net_73637;
  wire net_73643;
  wire net_73649;
  wire net_73653;
  wire net_73654;
  wire net_73697;
  wire net_73698;
  wire net_73700;
  wire net_73701;
  wire net_73702;
  wire net_73703;
  wire net_73704;
  wire net_73705;
  wire net_73706;
  wire net_73707;
  wire net_73708;
  wire net_73709;
  wire net_73711;
  wire net_73722;
  wire net_73723;
  wire net_73724;
  wire net_73728;
  wire net_73730;
  wire net_73731;
  wire net_73734;
  wire net_73736;
  wire net_73737;
  wire net_73738;
  wire net_73740;
  wire net_73742;
  wire net_73743;
  wire net_73744;
  wire net_73746;
  wire net_73748;
  wire net_73749;
  wire net_73750;
  wire net_73752;
  wire net_73754;
  wire net_73755;
  wire net_73756;
  wire net_73758;
  wire net_73760;
  wire net_73761;
  wire net_73762;
  wire net_73764;
  wire net_73766;
  wire net_73767;
  wire net_73768;
  wire net_73770;
  wire net_73772;
  wire net_73773;
  wire net_73774;
  wire net_73814;
  wire net_73819;
  wire net_73830;
  wire net_73835;
  wire net_73839;
  wire net_73841;
  wire net_73843;
  wire net_73844;
  wire net_73848;
  wire net_73850;
  wire net_73852;
  wire net_73853;
  wire net_73854;
  wire net_73855;
  wire net_73859;
  wire net_73864;
  wire net_73876;
  wire net_73878;
  wire net_73883;
  wire net_73895;
  wire net_73899;
  wire net_73900;
  wire net_73973;
  wire net_73999;
  wire net_74022;
  wire net_74023;
  wire net_75668;
  wire net_75671;
  wire net_75679;
  wire net_75682;
  wire net_75801;
  wire net_75806;
  wire net_75937;
  wire net_75938;
  wire net_75940;
  wire net_75942;
  wire net_75943;
  wire net_75944;
  wire net_76040;
  wire net_76141;
  wire net_76142;
  wire net_76143;
  wire net_76144;
  wire net_76145;
  wire net_76146;
  wire net_76147;
  wire net_76148;
  wire net_76192;
  wire net_76243;
  wire net_76247;
  wire net_76248;
  wire net_76290;
  wire net_76292;
  wire net_76300;
  wire net_76350;
  wire net_76453;
  wire net_76506;
  wire net_76511;
  wire net_76552;
  wire net_76553;
  wire net_76554;
  wire net_76556;
  wire net_76592;
  wire net_76651;
  wire net_76652;
  wire net_76655;
  wire net_76656;
  wire net_76710;
  wire net_76759;
  wire net_76760;
  wire net_76857;
  wire net_77062;
  wire net_79130;
  wire net_79143;
  wire net_79155;
  wire net_79173;
  wire net_79175;
  wire net_79204;
  wire net_79206;
  wire net_79207;
  wire net_79208;
  wire net_79209;
  wire net_79210;
  wire net_79212;
  wire net_79213;
  wire net_79217;
  wire net_79241;
  wire net_79259;
  wire net_79260;
  wire net_79268;
  wire net_79270;
  wire net_79278;
  wire net_79279;
  wire net_79287;
  wire net_79293;
  wire net_79302;
  wire net_79314;
  wire net_79320;
  wire net_79326;
  wire net_79331;
  wire net_79332;
  wire net_79333;
  wire net_79334;
  wire net_79335;
  wire net_79338;
  wire net_79340;
  wire net_79387;
  wire net_79388;
  wire net_79401;
  wire net_79414;
  wire net_79415;
  wire net_79453;
  wire net_79454;
  wire net_79455;
  wire net_79458;
  wire net_79460;
  wire net_79462;
  wire net_79475;
  wire net_79477;
  wire net_79501;
  wire net_79504;
  wire net_79505;
  wire net_79508;
  wire net_79519;
  wire net_79522;
  wire net_79527;
  wire net_79528;
  wire net_79530;
  wire net_79538;
  wire net_79543;
  wire net_79551;
  wire net_79554;
  wire net_79563;
  wire net_79569;
  wire net_79573;
  wire net_79577;
  wire net_79578;
  wire net_79583;
  wire net_79584;
  wire net_79585;
  wire net_79586;
  wire net_79595;
  wire net_79598;
  wire net_79601;
  wire net_79630;
  wire net_79631;
  wire net_79632;
  wire net_79633;
  wire net_79640;
  wire net_79641;
  wire net_79642;
  wire net_79645;
  wire net_79646;
  wire net_79647;
  wire net_79649;
  wire net_79653;
  wire net_79654;
  wire net_79655;
  wire net_79656;
  wire net_79677;
  wire net_79678;
  wire net_79679;
  wire net_79680;
  wire net_79683;
  wire net_79684;
  wire net_79685;
  wire net_79686;
  wire net_79699;
  wire net_79700;
  wire net_79701;
  wire net_79703;
  wire net_79704;
  wire net_79705;
  wire net_79709;
  wire net_79719;
  wire net_79745;
  wire net_79750;
  wire net_79752;
  wire net_79757;
  wire net_79770;
  wire net_79806;
  wire net_79807;
  wire net_79808;
  wire net_79809;
  wire net_79822;
  wire net_79823;
  wire net_79824;
  wire net_79826;
  wire net_79827;
  wire net_79828;
  wire net_79829;
  wire net_79830;
  wire net_79831;
  wire net_79832;
  wire net_79852;
  wire net_79855;
  wire net_79893;
  wire net_79937;
  wire net_79946;
  wire net_79947;
  wire net_79948;
  wire net_79949;
  wire net_79950;
  wire net_79951;
  wire net_79952;
  wire net_79954;
  wire net_79955;
  wire net_79996;
  wire net_79998;
  wire net_80004;
  wire net_80020;
  wire net_80043;
  wire net_80048;
  wire net_80053;
  wire net_80066;
  wire net_80069;
  wire net_80070;
  wire net_80071;
  wire net_80072;
  wire net_80073;
  wire net_80074;
  wire net_80075;
  wire net_80088;
  wire net_80093;
  wire net_80094;
  wire net_80113;
  wire net_80114;
  wire net_80118;
  wire net_80119;
  wire net_80126;
  wire net_80127;
  wire net_80146;
  wire net_80148;
  wire net_80151;
  wire net_80152;
  wire net_80169;
  wire net_80170;
  wire net_80175;
  wire net_80177;
  wire net_80191;
  wire net_80192;
  wire net_80193;
  wire net_80216;
  wire net_80242;
  wire net_80244;
  wire net_80307;
  wire net_80311;
  wire net_80315;
  wire net_80316;
  wire net_80362;
  wire net_80383;
  wire net_80403;
  wire net_80405;
  wire net_80437;
  wire net_80438;
  wire net_80439;
  wire net_80615;
  wire net_80631;
  wire net_80658;
  wire net_80683;
  wire net_80684;
  wire net_82732;
  wire net_82750;
  wire net_83041;
  wire net_83043;
  wire net_83045;
  wire net_83100;
  wire net_83102;
  wire net_83106;
  wire net_83112;
  wire net_83115;
  wire net_83130;
  wire net_83134;
  wire net_83157;
  wire net_83162;
  wire net_83163;
  wire net_83166;
  wire net_83170;
  wire net_83171;
  wire net_83176;
  wire net_83206;
  wire net_83219;
  wire net_83227;
  wire net_83228;
  wire net_83236;
  wire net_83238;
  wire net_83244;
  wire net_83252;
  wire net_83270;
  wire net_83280;
  wire net_83285;
  wire net_83286;
  wire net_83287;
  wire net_83290;
  wire net_83291;
  wire net_83293;
  wire net_83294;
  wire net_83328;
  wire net_83356;
  wire net_83357;
  wire net_83376;
  wire net_83385;
  wire net_83399;
  wire net_83408;
  wire net_83409;
  wire net_83414;
  wire net_83416;
  wire net_83427;
  wire net_83452;
  wire net_83471;
  wire net_83479;
  wire net_83481;
  wire net_83509;
  wire net_83514;
  wire net_83522;
  wire net_83526;
  wire net_83531;
  wire net_83532;
  wire net_83535;
  wire net_83537;
  wire net_83538;
  wire net_83540;
  wire net_83546;
  wire net_83576;
  wire net_83577;
  wire net_83579;
  wire net_83600;
  wire net_83614;
  wire net_83622;
  wire net_83627;
  wire net_83649;
  wire net_83654;
  wire net_83655;
  wire net_83656;
  wire net_83658;
  wire net_83659;
  wire net_83660;
  wire net_83661;
  wire net_83662;
  wire net_83681;
  wire net_83699;
  wire net_83701;
  wire net_83703;
  wire net_83704;
  wire net_83706;
  wire net_83707;
  wire net_83710;
  wire net_83711;
  wire net_83716;
  wire net_83717;
  wire net_83719;
  wire net_83720;
  wire net_83721;
  wire net_83725;
  wire net_83726;
  wire net_83727;
  wire net_83729;
  wire net_83731;
  wire net_83732;
  wire net_83735;
  wire net_83737;
  wire net_83738;
  wire net_83739;
  wire net_83741;
  wire net_83743;
  wire net_83744;
  wire net_83745;
  wire net_83747;
  wire net_83749;
  wire net_83750;
  wire net_83751;
  wire net_83753;
  wire net_83755;
  wire net_83756;
  wire net_83757;
  wire net_83759;
  wire net_83761;
  wire net_83762;
  wire net_83763;
  wire net_83765;
  wire net_83767;
  wire net_83768;
  wire net_83769;
  wire net_83771;
  wire net_83773;
  wire net_83774;
  wire net_83775;
  wire net_83777;
  wire net_83778;
  wire net_83779;
  wire net_83782;
  wire net_83783;
  wire net_83785;
  wire net_83786;
  wire net_83799;
  wire net_83815;
  wire net_83825;
  wire net_83830;
  wire net_83831;
  wire net_83832;
  wire net_83834;
  wire net_83835;
  wire net_83836;
  wire net_83840;
  wire net_83847;
  wire net_83850;
  wire net_83852;
  wire net_83854;
  wire net_83855;
  wire net_83856;
  wire net_83858;
  wire net_83860;
  wire net_83861;
  wire net_83862;
  wire net_83864;
  wire net_83866;
  wire net_83867;
  wire net_83868;
  wire net_83874;
  wire net_83877;
  wire net_83889;
  wire net_83895;
  wire net_83897;
  wire net_83900;
  wire net_83901;
  wire net_83902;
  wire net_83935;
  wire net_83943;
  wire net_83951;
  wire net_83954;
  wire net_83956;
  wire net_83958;
  wire net_83976;
  wire net_83983;
  wire net_83990;
  wire net_83995;
  wire net_84001;
  wire net_84023;
  wire net_84024;
  wire net_84037;
  wire net_84041;
  wire net_86563;
  wire net_86583;
  wire net_86709;
  wire net_86737;
  wire net_86745;
  wire net_86917;
  wire net_86924;
  wire net_86940;
  wire net_86948;
  wire net_86960;
  wire net_86972;
  wire net_86993;
  wire net_86994;
  wire net_87017;
  wire net_87036;
  wire net_87054;
  wire net_87059;
  wire net_87083;
  wire net_87105;
  wire net_87113;
  wire net_87116;
  wire net_87117;
  wire net_87118;
  wire net_87119;
  wire net_87122;
  wire net_87123;
  wire net_87125;
  wire net_87145;
  wire net_87163;
  wire net_87176;
  wire net_87177;
  wire net_87178;
  wire net_87183;
  wire net_87192;
  wire net_87210;
  wire net_87218;
  wire net_87231;
  wire net_87236;
  wire net_87239;
  wire net_87240;
  wire net_87242;
  wire net_87244;
  wire net_87248;
  wire net_87254;
  wire net_87256;
  wire net_87258;
  wire net_87262;
  wire net_87264;
  wire net_87301;
  wire net_87305;
  wire net_87342;
  wire net_87354;
  wire net_87362;
  wire net_87363;
  wire net_87375;
  wire net_87377;
  wire net_87383;
  wire net_87413;
  wire net_87428;
  wire net_87430;
  wire net_87434;
  wire net_87453;
  wire net_87465;
  wire net_87469;
  wire net_87483;
  wire net_87485;
  wire net_87486;
  wire net_87494;
  wire net_87502;
  wire net_87508;
  wire net_87510;
  wire net_87539;
  wire net_87542;
  wire net_87543;
  wire net_87547;
  wire net_87550;
  wire net_87557;
  wire net_87563;
  wire net_87575;
  wire net_87582;
  wire net_87588;
  wire net_87594;
  wire net_87600;
  wire net_87608;
  wire net_87609;
  wire net_87613;
  wire net_87629;
  wire net_87631;
  wire net_87633;
  wire net_87639;
  wire net_87665;
  wire net_87668;
  wire net_87676;
  wire net_87677;
  wire net_87682;
  wire net_87684;
  wire net_87702;
  wire net_87709;
  wire net_87721;
  wire net_87727;
  wire net_87731;
  wire net_87732;
  wire net_87765;
  wire net_87869;
  wire net_87871;
  wire net_87873;
  wire net_87992;
  wire net_87994;
  wire net_88117;
  wire net_88121;
  wire net_88242;
  wire net_88244;
  wire net_88248;
  wire net_90394;
  wire net_90410;
  wire net_90991;
  wire net_91009;
  wire net_91014;
  wire net_91018;
  wire net_91021;
  wire net_91023;
  wire net_91031;
  wire net_91048;
  wire net_91053;
  wire net_91067;
  wire net_91070;
  wire net_91071;
  wire net_91084;
  wire net_91094;
  wire net_91133;
  wire net_91137;
  wire net_91141;
  wire net_91152;
  wire net_91165;
  wire net_91188;
  wire net_91193;
  wire net_91194;
  wire net_91209;
  wire net_91217;
  wire net_91330;
  wire net_91380;
  wire net_91434;
  wire net_91439;
  wire net_91440;
  wire net_91463;
  wire net_91495;
  wire net_91536;
  wire net_91562;
  wire net_91563;
  wire net_91699;
  wire net_91701;
  wire net_91703;
  wire net_91705;
  wire net_91951;
  wire net_92076;
  wire net_94841;
  wire net_94843;
  wire net_94851;
  wire net_94984;
  wire net_94986;
  wire net_94987;
  wire net_95107;
  wire net_95109;
  wire net_95124;
  wire net_95128;
  wire net_95258;
  wire net_95259;
  wire net_95264;
  wire net_95397;
  wire net_95405;
  wire net_95407;
  wire net_95535;
  wire net_95538;
  wire net_95542;
  wire net_95545;
  wire net_95546;
  wire net_95675;
  wire net_95677;
  wire net_95678;
  wire net_95682;
  wire net_95685;
  wire net_96090;
  wire net_99270;
  wire net_99271;
  wire net_99272;
  wire net_99273;
  wire net_99274;
  wire net_99275;
  wire net_99276;
  wire net_99277;
  wire net_99370;
  wire net_99373;
  wire net_99380;
  wire net_99383;
  wire net_99385;
  wire net_99386;
  wire net_99388;
  wire net_99389;
  wire net_99391;
  wire net_99394;
  wire net_99395;
  wire net_99396;
  wire net_99398;
  wire net_99399;
  wire net_99400;
  wire net_99401;
  wire net_99403;
  wire net_99404;
  wire net_99405;
  wire net_99406;
  wire net_99407;
  wire net_99408;
  wire net_99409;
  wire net_99410;
  wire net_99411;
  wire net_99412;
  wire net_99413;
  wire net_99414;
  wire net_99415;
  wire net_99416;
  wire net_99417;
  wire net_99418;
  wire net_99420;
  wire net_99421;
  wire net_99422;
  wire net_99423;
  wire net_99424;
  wire net_99425;
  wire net_99426;
  wire net_99427;
  wire net_99458;
  wire net_99520;
  wire net_99521;
  wire net_99523;
  wire net_99527;
  wire net_99529;
  wire net_99530;
  wire net_99532;
  wire net_99533;
  wire net_99534;
  wire net_99535;
  wire net_99536;
  wire net_99543;
  wire net_99544;
  wire net_99545;
  wire net_99547;
  wire net_99549;
  wire net_99553;
  wire net_99554;
  wire net_99555;
  wire net_99556;
  wire net_99557;
  wire net_99558;
  wire net_99559;
  wire net_99560;
  wire net_99561;
  wire net_99562;
  wire net_99563;
  wire net_99564;
  wire net_99565;
  wire net_99566;
  wire net_99567;
  wire net_99568;
  wire net_99572;
  wire net_99573;
  wire net_99574;
  wire net_99575;
  wire net_99576;
  wire net_99577;
  wire net_99578;
  wire net_99579;
  wire net_99724;
  wire net_99725;
  wire net_99726;
  wire net_99727;
  wire net_99728;
  wire net_99729;
  wire net_99730;
  wire net_99731;
  wire net_100050;
  wire net_100051;
  wire net_100052;
  wire net_100053;
  wire net_100054;
  wire net_100055;
  wire net_100056;
  wire net_100057;
  wire net_100150;
  wire net_100154;
  wire net_100155;
  wire net_100156;
  wire net_100164;
  wire net_100168;
  wire net_100169;
  wire net_100170;
  wire net_100171;
  wire net_100172;
  wire net_100173;
  wire net_100175;
  wire net_100176;
  wire net_100178;
  wire net_100180;
  wire net_100181;
  wire net_100183;
  wire net_100184;
  wire net_100185;
  wire net_100186;
  wire net_100187;
  wire net_100188;
  wire net_100189;
  wire net_100190;
  wire net_100191;
  wire net_100192;
  wire net_100193;
  wire net_100194;
  wire net_100195;
  wire net_100196;
  wire net_100197;
  wire net_100198;
  wire net_100200;
  wire net_100201;
  wire net_100202;
  wire net_100203;
  wire net_100204;
  wire net_100205;
  wire net_100206;
  wire net_100207;
  wire net_100240;
  wire net_100302;
  wire net_100303;
  wire net_100309;
  wire net_100310;
  wire net_100311;
  wire net_100312;
  wire net_100313;
  wire net_100314;
  wire net_100317;
  wire net_100318;
  wire net_100319;
  wire net_100320;
  wire net_100325;
  wire net_100326;
  wire net_100330;
  wire net_100331;
  wire net_100333;
  wire net_100334;
  wire net_100335;
  wire net_100336;
  wire net_100337;
  wire net_100338;
  wire net_100339;
  wire net_100340;
  wire net_100341;
  wire net_100342;
  wire net_100343;
  wire net_100344;
  wire net_100345;
  wire net_100346;
  wire net_100347;
  wire net_100348;
  wire net_100352;
  wire net_100353;
  wire net_100354;
  wire net_100355;
  wire net_100356;
  wire net_100357;
  wire net_100358;
  wire net_100359;
  wire net_100504;
  wire net_100505;
  wire net_100506;
  wire net_100507;
  wire net_100508;
  wire net_100509;
  wire net_100510;
  wire net_100511;
  wire dangling_wire_0;
  wire dangling_wire_1;
  wire dangling_wire_10;
  wire dangling_wire_100;
  wire dangling_wire_101;
  wire dangling_wire_102;
  wire dangling_wire_103;
  wire dangling_wire_104;
  wire dangling_wire_105;
  wire dangling_wire_106;
  wire dangling_wire_107;
  wire dangling_wire_108;
  wire dangling_wire_109;
  wire dangling_wire_11;
  wire dangling_wire_110;
  wire dangling_wire_111;
  wire dangling_wire_112;
  wire dangling_wire_113;
  wire dangling_wire_114;
  wire dangling_wire_115;
  wire dangling_wire_116;
  wire dangling_wire_117;
  wire dangling_wire_118;
  wire dangling_wire_119;
  wire dangling_wire_12;
  wire dangling_wire_120;
  wire dangling_wire_121;
  wire dangling_wire_122;
  wire dangling_wire_123;
  wire dangling_wire_124;
  wire dangling_wire_125;
  wire dangling_wire_13;
  wire dangling_wire_14;
  wire dangling_wire_15;
  wire dangling_wire_16;
  wire dangling_wire_17;
  wire dangling_wire_18;
  wire dangling_wire_19;
  wire dangling_wire_2;
  wire dangling_wire_20;
  wire dangling_wire_21;
  wire dangling_wire_22;
  wire dangling_wire_23;
  wire dangling_wire_24;
  wire dangling_wire_25;
  wire dangling_wire_26;
  wire dangling_wire_27;
  wire dangling_wire_28;
  wire dangling_wire_29;
  wire dangling_wire_3;
  wire dangling_wire_30;
  wire dangling_wire_31;
  wire dangling_wire_32;
  wire dangling_wire_33;
  wire dangling_wire_34;
  wire dangling_wire_35;
  wire dangling_wire_36;
  wire dangling_wire_37;
  wire dangling_wire_38;
  wire dangling_wire_39;
  wire dangling_wire_4;
  wire dangling_wire_40;
  wire dangling_wire_41;
  wire dangling_wire_42;
  wire dangling_wire_43;
  wire dangling_wire_44;
  wire dangling_wire_45;
  wire dangling_wire_46;
  wire dangling_wire_47;
  wire dangling_wire_48;
  wire dangling_wire_49;
  wire dangling_wire_5;
  wire dangling_wire_50;
  wire dangling_wire_51;
  wire dangling_wire_52;
  wire dangling_wire_53;
  wire dangling_wire_54;
  wire dangling_wire_55;
  wire dangling_wire_56;
  wire dangling_wire_57;
  wire dangling_wire_58;
  wire dangling_wire_59;
  wire dangling_wire_6;
  wire dangling_wire_60;
  wire dangling_wire_61;
  wire dangling_wire_62;
  wire dangling_wire_63;
  wire dangling_wire_64;
  wire dangling_wire_65;
  wire dangling_wire_66;
  wire dangling_wire_67;
  wire dangling_wire_68;
  wire dangling_wire_69;
  wire dangling_wire_7;
  wire dangling_wire_70;
  wire dangling_wire_71;
  wire dangling_wire_72;
  wire dangling_wire_73;
  wire dangling_wire_74;
  wire dangling_wire_75;
  wire dangling_wire_76;
  wire dangling_wire_77;
  wire dangling_wire_78;
  wire dangling_wire_79;
  wire dangling_wire_8;
  wire dangling_wire_80;
  wire dangling_wire_81;
  wire dangling_wire_82;
  wire dangling_wire_83;
  wire dangling_wire_84;
  wire dangling_wire_85;
  wire dangling_wire_86;
  wire dangling_wire_87;
  wire dangling_wire_88;
  wire dangling_wire_89;
  wire dangling_wire_9;
  wire dangling_wire_90;
  wire dangling_wire_91;
  wire dangling_wire_92;
  wire dangling_wire_93;
  wire dangling_wire_94;
  wire dangling_wire_95;
  wire dangling_wire_96;
  wire dangling_wire_97;
  wire dangling_wire_98;
  wire dangling_wire_99;
  wire net_11324_cascademuxed;
  wire net_11336_cascademuxed;
  wire net_11348_cascademuxed;
  wire net_11469_cascademuxed;
  wire net_11475_cascademuxed;
  wire net_11481_cascademuxed;
  wire net_11487_cascademuxed;
  wire net_11499_cascademuxed;
  wire net_11505_cascademuxed;
  wire net_11511_cascademuxed;
  wire net_11598_cascademuxed;
  wire net_11616_cascademuxed;
  wire net_11622_cascademuxed;
  wire net_11628_cascademuxed;
  wire net_11634_cascademuxed;
  wire net_11715_cascademuxed;
  wire net_11733_cascademuxed;
  wire net_11739_cascademuxed;
  wire net_11745_cascademuxed;
  wire net_11751_cascademuxed;
  wire net_11838_cascademuxed;
  wire net_11850_cascademuxed;
  wire net_11862_cascademuxed;
  wire net_11967_cascademuxed;
  wire net_11973_cascademuxed;
  wire net_11979_cascademuxed;
  wire net_11991_cascademuxed;
  wire net_12090_cascademuxed;
  wire net_12120_cascademuxed;
  wire net_12207_cascademuxed;
  wire net_12213_cascademuxed;
  wire net_12225_cascademuxed;
  wire net_12231_cascademuxed;
  wire net_12249_cascademuxed;
  wire net_12477_cascademuxed;
  wire net_12483_cascademuxed;
  wire net_12573;
  wire net_12576_cascademuxed;
  wire net_12579;
  wire net_12582_cascademuxed;
  wire net_12585;
  wire net_12588_cascademuxed;
  wire net_12591;
  wire net_12594_cascademuxed;
  wire net_12597;
  wire net_12600_cascademuxed;
  wire net_12603;
  wire net_12606_cascademuxed;
  wire net_12609;
  wire net_12612_cascademuxed;
  wire net_12618_cascademuxed;
  wire net_12696;
  wire net_12699_cascademuxed;
  wire net_12702;
  wire net_12705_cascademuxed;
  wire net_12708;
  wire net_12711_cascademuxed;
  wire net_12714;
  wire net_12717_cascademuxed;
  wire net_12720;
  wire net_12723_cascademuxed;
  wire net_12726;
  wire net_12729_cascademuxed;
  wire net_12732;
  wire net_12735_cascademuxed;
  wire net_12741_cascademuxed;
  wire net_12822_cascademuxed;
  wire net_12828_cascademuxed;
  wire net_12840_cascademuxed;
  wire net_12942;
  wire net_12945_cascademuxed;
  wire net_12951_cascademuxed;
  wire net_12957_cascademuxed;
  wire net_12975_cascademuxed;
  wire net_13065;
  wire net_13068_cascademuxed;
  wire net_13074_cascademuxed;
  wire net_13080_cascademuxed;
  wire net_13086_cascademuxed;
  wire net_13203_cascademuxed;
  wire net_13227_cascademuxed;
  wire net_13233_cascademuxed;
  wire net_13356_cascademuxed;
  wire net_13479_cascademuxed;
  wire net_13560_cascademuxed;
  wire net_13596_cascademuxed;
  wire net_13959_cascademuxed;
  wire net_15137_cascademuxed;
  wire net_15143_cascademuxed;
  wire net_15149_cascademuxed;
  wire net_15155_cascademuxed;
  wire net_15173_cascademuxed;
  wire net_15179_cascademuxed;
  wire net_15300_cascademuxed;
  wire net_15306_cascademuxed;
  wire net_15312_cascademuxed;
  wire net_15318_cascademuxed;
  wire net_15330_cascademuxed;
  wire net_15342_cascademuxed;
  wire net_15423_cascademuxed;
  wire net_15429_cascademuxed;
  wire net_15441_cascademuxed;
  wire net_15447_cascademuxed;
  wire net_15453_cascademuxed;
  wire net_15459_cascademuxed;
  wire net_15465_cascademuxed;
  wire net_15546_cascademuxed;
  wire net_15564_cascademuxed;
  wire net_15570_cascademuxed;
  wire net_15705_cascademuxed;
  wire net_15816_cascademuxed;
  wire net_15828_cascademuxed;
  wire net_15912;
  wire net_15915_cascademuxed;
  wire net_15918;
  wire net_15921_cascademuxed;
  wire net_15924;
  wire net_15927_cascademuxed;
  wire net_15930;
  wire net_15933_cascademuxed;
  wire net_15936;
  wire net_15939_cascademuxed;
  wire net_15942;
  wire net_15945_cascademuxed;
  wire net_15957_cascademuxed;
  wire net_16038_cascademuxed;
  wire net_16158;
  wire net_16161_cascademuxed;
  wire net_16164;
  wire net_16167_cascademuxed;
  wire net_16170;
  wire net_16173_cascademuxed;
  wire net_16176;
  wire net_16179_cascademuxed;
  wire net_16182;
  wire net_16185_cascademuxed;
  wire net_16188;
  wire net_16191_cascademuxed;
  wire net_16197_cascademuxed;
  wire net_16296_cascademuxed;
  wire net_16320_cascademuxed;
  wire net_16326_cascademuxed;
  wire net_16419_cascademuxed;
  wire net_16425_cascademuxed;
  wire net_16431_cascademuxed;
  wire net_16443_cascademuxed;
  wire net_16527;
  wire net_16530_cascademuxed;
  wire net_16533;
  wire net_16536_cascademuxed;
  wire net_16539;
  wire net_16542_cascademuxed;
  wire net_16545;
  wire net_16548_cascademuxed;
  wire net_16551;
  wire net_16554_cascademuxed;
  wire net_16557;
  wire net_16560_cascademuxed;
  wire net_16566_cascademuxed;
  wire net_16650;
  wire net_16653_cascademuxed;
  wire net_16656;
  wire net_16659_cascademuxed;
  wire net_16662;
  wire net_16665_cascademuxed;
  wire net_16668;
  wire net_16671_cascademuxed;
  wire net_16674;
  wire net_16677_cascademuxed;
  wire net_16680;
  wire net_16683_cascademuxed;
  wire net_16686;
  wire net_16689_cascademuxed;
  wire net_16695_cascademuxed;
  wire net_16776_cascademuxed;
  wire net_16782_cascademuxed;
  wire net_16794_cascademuxed;
  wire net_16812_cascademuxed;
  wire net_16896;
  wire net_16899_cascademuxed;
  wire net_16902;
  wire net_16905_cascademuxed;
  wire net_16908;
  wire net_16911_cascademuxed;
  wire net_16914;
  wire net_16917_cascademuxed;
  wire net_16920;
  wire net_16923_cascademuxed;
  wire net_16926;
  wire net_16929_cascademuxed;
  wire net_16935_cascademuxed;
  wire net_17169_cascademuxed;
  wire net_17268_cascademuxed;
  wire net_17298_cascademuxed;
  wire net_17304_cascademuxed;
  wire net_17421_cascademuxed;
  wire net_18968_cascademuxed;
  wire net_18980_cascademuxed;
  wire net_18992_cascademuxed;
  wire net_18998_cascademuxed;
  wire net_19004_cascademuxed;
  wire net_19010_cascademuxed;
  wire net_19128;
  wire net_19131_cascademuxed;
  wire net_19134;
  wire net_19137_cascademuxed;
  wire net_19140;
  wire net_19143_cascademuxed;
  wire net_19146;
  wire net_19149_cascademuxed;
  wire net_19152;
  wire net_19155_cascademuxed;
  wire net_19158;
  wire net_19161_cascademuxed;
  wire net_19164;
  wire net_19167_cascademuxed;
  wire net_19173_cascademuxed;
  wire net_19251;
  wire net_19254_cascademuxed;
  wire net_19257;
  wire net_19260_cascademuxed;
  wire net_19263;
  wire net_19266_cascademuxed;
  wire net_19272_cascademuxed;
  wire net_19284_cascademuxed;
  wire net_19290_cascademuxed;
  wire net_19296_cascademuxed;
  wire net_19377_cascademuxed;
  wire net_19395_cascademuxed;
  wire net_19401_cascademuxed;
  wire net_19413_cascademuxed;
  wire net_19500_cascademuxed;
  wire net_19524_cascademuxed;
  wire net_19530_cascademuxed;
  wire net_19536_cascademuxed;
  wire net_19623_cascademuxed;
  wire net_19629_cascademuxed;
  wire net_19641_cascademuxed;
  wire net_19647_cascademuxed;
  wire net_19653_cascademuxed;
  wire net_19659_cascademuxed;
  wire net_19746_cascademuxed;
  wire net_19758_cascademuxed;
  wire net_19764_cascademuxed;
  wire net_19770_cascademuxed;
  wire net_19788_cascademuxed;
  wire net_19869_cascademuxed;
  wire net_19875_cascademuxed;
  wire net_19881_cascademuxed;
  wire net_19887_cascademuxed;
  wire net_19893_cascademuxed;
  wire net_19899_cascademuxed;
  wire net_19902;
  wire net_19905_cascademuxed;
  wire net_19911_cascademuxed;
  wire net_19989;
  wire net_19992_cascademuxed;
  wire net_19995;
  wire net_19998_cascademuxed;
  wire net_20001;
  wire net_20004_cascademuxed;
  wire net_20007;
  wire net_20010_cascademuxed;
  wire net_20013;
  wire net_20016_cascademuxed;
  wire net_20019;
  wire net_20022_cascademuxed;
  wire net_20025;
  wire net_20028_cascademuxed;
  wire net_20034_cascademuxed;
  wire net_20112;
  wire net_20115_cascademuxed;
  wire net_20118;
  wire net_20121_cascademuxed;
  wire net_20124;
  wire net_20127_cascademuxed;
  wire net_20130;
  wire net_20133_cascademuxed;
  wire net_20136;
  wire net_20139_cascademuxed;
  wire net_20142;
  wire net_20145_cascademuxed;
  wire net_20151_cascademuxed;
  wire net_20262_cascademuxed;
  wire net_20274_cascademuxed;
  wire net_20367_cascademuxed;
  wire net_20391_cascademuxed;
  wire net_20484_cascademuxed;
  wire net_20490_cascademuxed;
  wire net_20496_cascademuxed;
  wire net_20502_cascademuxed;
  wire net_20508_cascademuxed;
  wire net_20514_cascademuxed;
  wire net_20517;
  wire net_20520_cascademuxed;
  wire net_20625_cascademuxed;
  wire net_20637_cascademuxed;
  wire net_20766_cascademuxed;
  wire net_20877_cascademuxed;
  wire net_20883_cascademuxed;
  wire net_21006_cascademuxed;
  wire net_21117_cascademuxed;
  wire net_21222_cascademuxed;
  wire net_21258_cascademuxed;
  wire net_21264_cascademuxed;
  wire net_21375_cascademuxed;
  wire net_22817_cascademuxed;
  wire net_22841_cascademuxed;
  wire net_22968_cascademuxed;
  wire net_23127_cascademuxed;
  wire net_23220_cascademuxed;
  wire net_23232_cascademuxed;
  wire net_23328;
  wire net_23331_cascademuxed;
  wire net_23334;
  wire net_23340;
  wire net_23346;
  wire net_23352;
  wire net_23358;
  wire net_23361_cascademuxed;
  wire net_23364;
  wire net_23451;
  wire net_23454_cascademuxed;
  wire net_23457;
  wire net_23460_cascademuxed;
  wire net_23463;
  wire net_23466_cascademuxed;
  wire net_23469;
  wire net_23472_cascademuxed;
  wire net_23475;
  wire net_23478_cascademuxed;
  wire net_23481;
  wire net_23484_cascademuxed;
  wire net_23496_cascademuxed;
  wire net_23583_cascademuxed;
  wire net_23589_cascademuxed;
  wire net_23595_cascademuxed;
  wire net_23607_cascademuxed;
  wire net_23700_cascademuxed;
  wire net_23706_cascademuxed;
  wire net_23736_cascademuxed;
  wire net_23964_cascademuxed;
  wire net_24081_cascademuxed;
  wire net_24087_cascademuxed;
  wire net_24216_cascademuxed;
  wire net_24333_cascademuxed;
  wire net_24438_cascademuxed;
  wire net_24462_cascademuxed;
  wire net_24696_cascademuxed;
  wire net_24714_cascademuxed;
  wire net_24720_cascademuxed;
  wire net_24726_cascademuxed;
  wire net_24813_cascademuxed;
  wire net_24948_cascademuxed;
  wire net_25053_cascademuxed;
  wire net_25077_cascademuxed;
  wire net_26885_cascademuxed;
  wire net_26886_cascademuxed;
  wire net_26888_cascademuxed;
  wire net_26889_cascademuxed;
  wire net_26890_cascademuxed;
  wire net_26891_cascademuxed;
  wire net_26987_cascademuxed;
  wire net_26988_cascademuxed;
  wire net_26990_cascademuxed;
  wire net_26991_cascademuxed;
  wire net_26992_cascademuxed;
  wire net_26993_cascademuxed;
  wire net_27497_cascademuxed;
  wire net_27498_cascademuxed;
  wire net_27701_cascademuxed;
  wire net_27702_cascademuxed;
  wire net_30116_cascademuxed;
  wire net_30269_cascademuxed;
  wire net_30281_cascademuxed;
  wire net_30359;
  wire net_30362_cascademuxed;
  wire net_30365;
  wire net_30368_cascademuxed;
  wire net_30374_cascademuxed;
  wire net_30380_cascademuxed;
  wire net_30386_cascademuxed;
  wire net_30392_cascademuxed;
  wire net_30398_cascademuxed;
  wire net_30482;
  wire net_30485_cascademuxed;
  wire net_30488;
  wire net_30491_cascademuxed;
  wire net_30497_cascademuxed;
  wire net_30521_cascademuxed;
  wire net_30608_cascademuxed;
  wire net_30614_cascademuxed;
  wire net_30632_cascademuxed;
  wire net_30743_cascademuxed;
  wire net_30755_cascademuxed;
  wire net_30896_cascademuxed;
  wire net_30983_cascademuxed;
  wire net_31001_cascademuxed;
  wire net_31100_cascademuxed;
  wire net_31220;
  wire net_31223_cascademuxed;
  wire net_31226;
  wire net_31229_cascademuxed;
  wire net_31232;
  wire net_31235_cascademuxed;
  wire net_31238;
  wire net_31241_cascademuxed;
  wire net_31244;
  wire net_31247_cascademuxed;
  wire net_31250;
  wire net_31253_cascademuxed;
  wire net_31256;
  wire net_31259_cascademuxed;
  wire net_31364_cascademuxed;
  wire net_31376_cascademuxed;
  wire net_31382_cascademuxed;
  wire net_31505_cascademuxed;
  wire net_31511_cascademuxed;
  wire net_31592_cascademuxed;
  wire net_31598_cascademuxed;
  wire net_31604_cascademuxed;
  wire net_31610_cascademuxed;
  wire net_31616_cascademuxed;
  wire net_31622_cascademuxed;
  wire net_31628_cascademuxed;
  wire net_31634_cascademuxed;
  wire net_31727_cascademuxed;
  wire net_31838_cascademuxed;
  wire net_31844_cascademuxed;
  wire net_31850_cascademuxed;
  wire net_31856_cascademuxed;
  wire net_31862_cascademuxed;
  wire net_31868_cascademuxed;
  wire net_31874_cascademuxed;
  wire net_31961_cascademuxed;
  wire net_31979_cascademuxed;
  wire net_31991_cascademuxed;
  wire net_32084_cascademuxed;
  wire net_32102_cascademuxed;
  wire net_33673_cascademuxed;
  wire net_33824_cascademuxed;
  wire net_33947_cascademuxed;
  wire net_33983_cascademuxed;
  wire net_34205_cascademuxed;
  wire net_34217_cascademuxed;
  wire net_34235_cascademuxed;
  wire net_34346_cascademuxed;
  wire net_34439_cascademuxed;
  wire net_34559;
  wire net_34562_cascademuxed;
  wire net_34565;
  wire net_34568_cascademuxed;
  wire net_34571;
  wire net_34574_cascademuxed;
  wire net_34577;
  wire net_34580_cascademuxed;
  wire net_34583;
  wire net_34586_cascademuxed;
  wire net_34589;
  wire net_34592_cascademuxed;
  wire net_34595;
  wire net_34598_cascademuxed;
  wire net_34691_cascademuxed;
  wire net_34709_cascademuxed;
  wire net_34820_cascademuxed;
  wire net_34937_cascademuxed;
  wire net_35054_cascademuxed;
  wire net_35066_cascademuxed;
  wire net_35078_cascademuxed;
  wire net_35087;
  wire net_35189_cascademuxed;
  wire net_35207_cascademuxed;
  wire net_35336_cascademuxed;
  wire net_35423_cascademuxed;
  wire net_35429_cascademuxed;
  wire net_35435_cascademuxed;
  wire net_35441_cascademuxed;
  wire net_35447_cascademuxed;
  wire net_35459_cascademuxed;
  wire net_35465_cascademuxed;
  wire net_35552_cascademuxed;
  wire net_35564_cascademuxed;
  wire net_35582_cascademuxed;
  wire net_37498_cascademuxed;
  wire net_37510_cascademuxed;
  wire net_37516_cascademuxed;
  wire net_37691_cascademuxed;
  wire net_37814_cascademuxed;
  wire net_37901_cascademuxed;
  wire net_37937_cascademuxed;
  wire net_38024_cascademuxed;
  wire net_38060_cascademuxed;
  wire net_38276_cascademuxed;
  wire net_38294_cascademuxed;
  wire net_38312_cascademuxed;
  wire net_38390;
  wire net_38393_cascademuxed;
  wire net_38396;
  wire net_38399_cascademuxed;
  wire net_38402;
  wire net_38408;
  wire net_38411_cascademuxed;
  wire net_38414;
  wire net_38420;
  wire net_38423_cascademuxed;
  wire net_38426;
  wire net_38429_cascademuxed;
  wire net_38435_cascademuxed;
  wire net_38522_cascademuxed;
  wire net_38528_cascademuxed;
  wire net_38639_cascademuxed;
  wire net_38675_cascademuxed;
  wire net_38891_cascademuxed;
  wire net_39026_cascademuxed;
  wire net_39044_cascademuxed;
  wire net_39131_cascademuxed;
  wire net_39254_cascademuxed;
  wire net_39260_cascademuxed;
  wire net_39266_cascademuxed;
  wire net_39272_cascademuxed;
  wire net_39278_cascademuxed;
  wire net_39284_cascademuxed;
  wire net_39401_cascademuxed;
  wire net_39419_cascademuxed;
  wire net_39506_cascademuxed;
  wire net_39512_cascademuxed;
  wire net_39518_cascademuxed;
  wire net_39623_cascademuxed;
  wire net_39629_cascademuxed;
  wire net_39635_cascademuxed;
  wire net_39653_cascademuxed;
  wire net_39659_cascademuxed;
  wire net_39665_cascademuxed;
  wire net_41320;
  wire net_41323_cascademuxed;
  wire net_41329_cascademuxed;
  wire net_41365_cascademuxed;
  wire net_41504_cascademuxed;
  wire net_41615_cascademuxed;
  wire net_41627_cascademuxed;
  wire net_41633_cascademuxed;
  wire net_41645_cascademuxed;
  wire net_41732_cascademuxed;
  wire net_41750_cascademuxed;
  wire net_41774_cascademuxed;
  wire net_42107_cascademuxed;
  wire net_42125_cascademuxed;
  wire net_42248_cascademuxed;
  wire net_42365_cascademuxed;
  wire net_42470_cascademuxed;
  wire net_42500_cascademuxed;
  wire net_42506_cascademuxed;
  wire net_42512_cascademuxed;
  wire net_42617_cascademuxed;
  wire net_42635_cascademuxed;
  wire net_42851_cascademuxed;
  wire net_42980_cascademuxed;
  wire net_43085_cascademuxed;
  wire net_43097_cascademuxed;
  wire net_43109_cascademuxed;
  wire net_43226_cascademuxed;
  wire net_43331_cascademuxed;
  wire net_43343_cascademuxed;
  wire net_43367_cascademuxed;
  wire net_43454_cascademuxed;
  wire net_43460_cascademuxed;
  wire net_43466_cascademuxed;
  wire net_43478_cascademuxed;
  wire net_43484_cascademuxed;
  wire net_43496_cascademuxed;
  wire net_43583_cascademuxed;
  wire net_43619_cascademuxed;
  wire net_45178_cascademuxed;
  wire net_45314;
  wire net_45317_cascademuxed;
  wire net_45323_cascademuxed;
  wire net_45329_cascademuxed;
  wire net_45347_cascademuxed;
  wire net_45353_cascademuxed;
  wire net_45437;
  wire net_45440_cascademuxed;
  wire net_45443;
  wire net_45446_cascademuxed;
  wire net_45449;
  wire net_45452_cascademuxed;
  wire net_45455;
  wire net_45458_cascademuxed;
  wire net_45461;
  wire net_45464_cascademuxed;
  wire net_45467;
  wire net_45470_cascademuxed;
  wire net_45473;
  wire net_45476_cascademuxed;
  wire net_45560;
  wire net_45563_cascademuxed;
  wire net_45566;
  wire net_45569_cascademuxed;
  wire net_45572;
  wire net_45575_cascademuxed;
  wire net_45578;
  wire net_45581_cascademuxed;
  wire net_45584;
  wire net_45587_cascademuxed;
  wire net_45590;
  wire net_45593_cascademuxed;
  wire net_45596;
  wire net_45599_cascademuxed;
  wire net_45605_cascademuxed;
  wire net_45692_cascademuxed;
  wire net_46055_cascademuxed;
  wire net_46061_cascademuxed;
  wire net_46079_cascademuxed;
  wire net_46307_cascademuxed;
  wire net_46343_cascademuxed;
  wire net_46424_cascademuxed;
  wire net_46442_cascademuxed;
  wire net_46547_cascademuxed;
  wire net_46553_cascademuxed;
  wire net_46571_cascademuxed;
  wire net_46577_cascademuxed;
  wire net_46682_cascademuxed;
  wire net_46694_cascademuxed;
  wire net_46817_cascademuxed;
  wire net_46928_cascademuxed;
  wire net_46958_cascademuxed;
  wire net_47039_cascademuxed;
  wire net_47045_cascademuxed;
  wire net_47057_cascademuxed;
  wire net_47063_cascademuxed;
  wire net_47162_cascademuxed;
  wire net_47192_cascademuxed;
  wire net_47198_cascademuxed;
  wire net_47291_cascademuxed;
  wire net_47297_cascademuxed;
  wire net_47315_cascademuxed;
  wire net_47327_cascademuxed;
  wire net_48985_cascademuxed;
  wire net_48988;
  wire net_48994;
  wire net_48997_cascademuxed;
  wire net_49009_cascademuxed;
  wire net_49148_cascademuxed;
  wire net_49271_cascademuxed;
  wire net_49289_cascademuxed;
  wire net_49295_cascademuxed;
  wire net_49400_cascademuxed;
  wire net_49418_cascademuxed;
  wire net_49430_cascademuxed;
  wire net_49517_cascademuxed;
  wire net_49640_cascademuxed;
  wire net_49670_cascademuxed;
  wire net_49763_cascademuxed;
  wire net_49781_cascademuxed;
  wire net_49886_cascademuxed;
  wire net_49916_cascademuxed;
  wire net_50168_cascademuxed;
  wire net_50174_cascademuxed;
  wire net_50279_cascademuxed;
  wire net_50285_cascademuxed;
  wire net_50291_cascademuxed;
  wire net_50396_cascademuxed;
  wire net_50501_cascademuxed;
  wire net_50624_cascademuxed;
  wire net_50630_cascademuxed;
  wire net_50642_cascademuxed;
  wire net_50648_cascademuxed;
  wire net_50654_cascademuxed;
  wire net_50753_cascademuxed;
  wire net_50759_cascademuxed;
  wire net_50765_cascademuxed;
  wire net_50771_cascademuxed;
  wire net_50777_cascademuxed;
  wire net_50789_cascademuxed;
  wire net_50870_cascademuxed;
  wire net_50876_cascademuxed;
  wire net_50882_cascademuxed;
  wire net_50888_cascademuxed;
  wire net_50894_cascademuxed;
  wire net_50900_cascademuxed;
  wire net_50906_cascademuxed;
  wire net_50912_cascademuxed;
  wire net_50993_cascademuxed;
  wire net_50999_cascademuxed;
  wire net_51011_cascademuxed;
  wire net_51035_cascademuxed;
  wire net_52846_cascademuxed;
  wire net_52852_cascademuxed;
  wire net_52985_cascademuxed;
  wire net_53126_cascademuxed;
  wire net_53132_cascademuxed;
  wire net_53138_cascademuxed;
  wire net_53144_cascademuxed;
  wire net_53231_cascademuxed;
  wire net_53261_cascademuxed;
  wire net_53354_cascademuxed;
  wire net_53384_cascademuxed;
  wire net_53495_cascademuxed;
  wire net_53600_cascademuxed;
  wire net_53606_cascademuxed;
  wire net_53624_cascademuxed;
  wire net_53630_cascademuxed;
  wire net_53636_cascademuxed;
  wire net_53717_cascademuxed;
  wire net_53723_cascademuxed;
  wire net_53729_cascademuxed;
  wire net_53741_cascademuxed;
  wire net_53747_cascademuxed;
  wire net_53753_cascademuxed;
  wire net_53852_cascademuxed;
  wire net_53963_cascademuxed;
  wire net_53969_cascademuxed;
  wire net_53987_cascademuxed;
  wire net_54110_cascademuxed;
  wire net_54116_cascademuxed;
  wire net_54122_cascademuxed;
  wire net_54245_cascademuxed;
  wire net_54251_cascademuxed;
  wire net_54338_cascademuxed;
  wire net_54356_cascademuxed;
  wire net_54368_cascademuxed;
  wire net_54374_cascademuxed;
  wire net_54461_cascademuxed;
  wire net_54491_cascademuxed;
  wire net_54497_cascademuxed;
  wire net_54578_cascademuxed;
  wire net_54584_cascademuxed;
  wire net_54590_cascademuxed;
  wire net_54620_cascademuxed;
  wire net_54707_cascademuxed;
  wire net_54719_cascademuxed;
  wire net_54725_cascademuxed;
  wire net_54731_cascademuxed;
  wire net_54737_cascademuxed;
  wire net_54842_cascademuxed;
  wire net_54854_cascademuxed;
  wire net_54947_cascademuxed;
  wire net_54953_cascademuxed;
  wire net_54959_cascademuxed;
  wire net_54965_cascademuxed;
  wire net_54977_cascademuxed;
  wire net_54983_cascademuxed;
  wire net_54989_cascademuxed;
  wire net_55112_cascademuxed;
  wire net_56682_cascademuxed;
  wire net_56809_cascademuxed;
  wire net_56827_cascademuxed;
  wire net_56845_cascademuxed;
  wire net_57055_cascademuxed;
  wire net_57067_cascademuxed;
  wire net_57079_cascademuxed;
  wire net_57178_cascademuxed;
  wire net_57202_cascademuxed;
  wire net_57208_cascademuxed;
  wire net_57214_cascademuxed;
  wire net_57307_cascademuxed;
  wire net_57319_cascademuxed;
  wire net_57325_cascademuxed;
  wire net_57337_cascademuxed;
  wire net_57343_cascademuxed;
  wire net_57460_cascademuxed;
  wire net_57547_cascademuxed;
  wire net_57559_cascademuxed;
  wire net_57583_cascademuxed;
  wire net_57706_cascademuxed;
  wire net_57799_cascademuxed;
  wire net_57817_cascademuxed;
  wire net_57835_cascademuxed;
  wire net_57934_cascademuxed;
  wire net_58174_cascademuxed;
  wire net_58180_cascademuxed;
  wire net_58186_cascademuxed;
  wire net_58198_cascademuxed;
  wire net_58204_cascademuxed;
  wire net_58285_cascademuxed;
  wire net_58321_cascademuxed;
  wire net_58327_cascademuxed;
  wire net_58444_cascademuxed;
  wire net_58531_cascademuxed;
  wire net_58534;
  wire net_58537_cascademuxed;
  wire net_58540;
  wire net_58543_cascademuxed;
  wire net_58546;
  wire net_58549_cascademuxed;
  wire net_58552;
  wire net_58555_cascademuxed;
  wire net_58558;
  wire net_58561_cascademuxed;
  wire net_58564;
  wire net_58567_cascademuxed;
  wire net_58573_cascademuxed;
  wire net_58654_cascademuxed;
  wire net_58672_cascademuxed;
  wire net_58690_cascademuxed;
  wire net_58777_cascademuxed;
  wire net_58783_cascademuxed;
  wire net_58789_cascademuxed;
  wire net_58795_cascademuxed;
  wire net_58807_cascademuxed;
  wire net_58813_cascademuxed;
  wire net_58819_cascademuxed;
  wire net_58918_cascademuxed;
  wire net_60774_cascademuxed;
  wire net_60909_cascademuxed;
  wire net_60915_cascademuxed;
  wire net_60921_cascademuxed;
  wire net_61020_cascademuxed;
  wire net_61032_cascademuxed;
  wire net_61044_cascademuxed;
  wire net_61131_cascademuxed;
  wire net_61137_cascademuxed;
  wire net_61149_cascademuxed;
  wire net_61155_cascademuxed;
  wire net_61161_cascademuxed;
  wire net_61167_cascademuxed;
  wire net_61173_cascademuxed;
  wire net_61266_cascademuxed;
  wire net_61272_cascademuxed;
  wire net_61290_cascademuxed;
  wire net_61395_cascademuxed;
  wire net_61506_cascademuxed;
  wire net_61524_cascademuxed;
  wire net_61536_cascademuxed;
  wire net_61626;
  wire net_61641_cascademuxed;
  wire net_61746_cascademuxed;
  wire net_61752_cascademuxed;
  wire net_61776_cascademuxed;
  wire net_61788_cascademuxed;
  wire net_61869_cascademuxed;
  wire net_61887_cascademuxed;
  wire net_61899_cascademuxed;
  wire net_61989;
  wire net_61992_cascademuxed;
  wire net_61995;
  wire net_62001;
  wire net_62004_cascademuxed;
  wire net_62007;
  wire net_62010_cascademuxed;
  wire net_62013;
  wire net_62019;
  wire net_62025;
  wire net_62115_cascademuxed;
  wire net_62121_cascademuxed;
  wire net_62127_cascademuxed;
  wire net_62133_cascademuxed;
  wire net_62145_cascademuxed;
  wire net_62250_cascademuxed;
  wire net_62256_cascademuxed;
  wire net_62280_cascademuxed;
  wire net_62361_cascademuxed;
  wire net_62364;
  wire net_62367_cascademuxed;
  wire net_62370;
  wire net_62373_cascademuxed;
  wire net_62376;
  wire net_62379_cascademuxed;
  wire net_62382;
  wire net_62385_cascademuxed;
  wire net_62388;
  wire net_62391_cascademuxed;
  wire net_62394;
  wire net_62397_cascademuxed;
  wire net_62403_cascademuxed;
  wire net_62481;
  wire net_62484_cascademuxed;
  wire net_62496_cascademuxed;
  wire net_62631_cascademuxed;
  wire net_64488_cascademuxed;
  wire net_64605_cascademuxed;
  wire net_64713;
  wire net_64716_cascademuxed;
  wire net_64719;
  wire net_64722_cascademuxed;
  wire net_64725;
  wire net_64728_cascademuxed;
  wire net_64731;
  wire net_64734_cascademuxed;
  wire net_64737;
  wire net_64740_cascademuxed;
  wire net_64743;
  wire net_64746_cascademuxed;
  wire net_64749;
  wire net_64752_cascademuxed;
  wire net_64758_cascademuxed;
  wire net_64836;
  wire net_64839_cascademuxed;
  wire net_64842;
  wire net_64845_cascademuxed;
  wire net_64848;
  wire net_64851_cascademuxed;
  wire net_64881_cascademuxed;
  wire net_64959;
  wire net_64962_cascademuxed;
  wire net_64965;
  wire net_64968_cascademuxed;
  wire net_64971;
  wire net_64974_cascademuxed;
  wire net_64977;
  wire net_64983;
  wire net_64986_cascademuxed;
  wire net_64989;
  wire net_64995;
  wire net_64998_cascademuxed;
  wire net_65004_cascademuxed;
  wire net_65082;
  wire net_65085_cascademuxed;
  wire net_65088;
  wire net_65094;
  wire net_65100;
  wire net_65103_cascademuxed;
  wire net_65121_cascademuxed;
  wire net_65214_cascademuxed;
  wire net_65232_cascademuxed;
  wire net_65337_cascademuxed;
  wire net_65454_cascademuxed;
  wire net_65472_cascademuxed;
  wire net_65478_cascademuxed;
  wire net_65574;
  wire net_65577_cascademuxed;
  wire net_65580;
  wire net_65583_cascademuxed;
  wire net_65586;
  wire net_65589_cascademuxed;
  wire net_65592;
  wire net_65595_cascademuxed;
  wire net_65598;
  wire net_65601_cascademuxed;
  wire net_65613_cascademuxed;
  wire net_65712_cascademuxed;
  wire net_65718_cascademuxed;
  wire net_65736_cascademuxed;
  wire net_65742_cascademuxed;
  wire net_65820;
  wire net_65823_cascademuxed;
  wire net_65826;
  wire net_65829_cascademuxed;
  wire net_65832;
  wire net_65835_cascademuxed;
  wire net_65838;
  wire net_65841_cascademuxed;
  wire net_65844;
  wire net_65847_cascademuxed;
  wire net_65850;
  wire net_65853_cascademuxed;
  wire net_65943;
  wire net_65946_cascademuxed;
  wire net_65949;
  wire net_65952_cascademuxed;
  wire net_65955;
  wire net_65958_cascademuxed;
  wire net_65961;
  wire net_65964_cascademuxed;
  wire net_65967;
  wire net_65970_cascademuxed;
  wire net_65973;
  wire net_65976_cascademuxed;
  wire net_65979;
  wire net_65982_cascademuxed;
  wire net_65988_cascademuxed;
  wire net_66069_cascademuxed;
  wire net_66075_cascademuxed;
  wire net_66105_cascademuxed;
  wire net_66192_cascademuxed;
  wire net_66198_cascademuxed;
  wire net_66204_cascademuxed;
  wire net_66210_cascademuxed;
  wire net_66216_cascademuxed;
  wire net_66228_cascademuxed;
  wire net_66234_cascademuxed;
  wire net_66315_cascademuxed;
  wire net_66321_cascademuxed;
  wire net_66327_cascademuxed;
  wire net_66345_cascademuxed;
  wire net_66357_cascademuxed;
  wire net_66438_cascademuxed;
  wire net_6792_cascademuxed;
  wire net_68424_cascademuxed;
  wire net_68430_cascademuxed;
  wire net_68436_cascademuxed;
  wire net_68553_cascademuxed;
  wire net_68583_cascademuxed;
  wire net_68589_cascademuxed;
  wire net_68670_cascademuxed;
  wire net_68682_cascademuxed;
  wire net_68706_cascademuxed;
  wire net_68712_cascademuxed;
  wire net_68805_cascademuxed;
  wire net_68835_cascademuxed;
  wire net_68958_cascademuxed;
  wire net_69045_cascademuxed;
  wire net_69051_cascademuxed;
  wire net_69075_cascademuxed;
  wire net_69303_cascademuxed;
  wire net_6937_cascademuxed;
  wire net_6940;
  wire net_69405;
  wire net_69408_cascademuxed;
  wire net_69411;
  wire net_69414_cascademuxed;
  wire net_69417;
  wire net_69420_cascademuxed;
  wire net_69423;
  wire net_69426_cascademuxed;
  wire net_69438_cascademuxed;
  wire net_6943_cascademuxed;
  wire net_6946;
  wire net_6949_cascademuxed;
  wire net_6952;
  wire net_69549_cascademuxed;
  wire net_69555_cascademuxed;
  wire net_6955_cascademuxed;
  wire net_6958;
  wire net_69651;
  wire net_69654_cascademuxed;
  wire net_69657;
  wire net_69660_cascademuxed;
  wire net_69663;
  wire net_69666_cascademuxed;
  wire net_69669;
  wire net_69672_cascademuxed;
  wire net_69675;
  wire net_69678_cascademuxed;
  wire net_6967_cascademuxed;
  wire net_69681;
  wire net_69684_cascademuxed;
  wire net_69690_cascademuxed;
  wire net_69696_cascademuxed;
  wire net_69777_cascademuxed;
  wire net_69783_cascademuxed;
  wire net_69789_cascademuxed;
  wire net_69795_cascademuxed;
  wire net_6979_cascademuxed;
  wire net_69801_cascademuxed;
  wire net_69813_cascademuxed;
  wire net_69819_cascademuxed;
  wire net_69900_cascademuxed;
  wire net_69918_cascademuxed;
  wire net_69930_cascademuxed;
  wire net_70020;
  wire net_70023_cascademuxed;
  wire net_70026;
  wire net_70032;
  wire net_70035_cascademuxed;
  wire net_70038;
  wire net_70041_cascademuxed;
  wire net_70044;
  wire net_70050;
  wire net_70152_cascademuxed;
  wire net_70170_cascademuxed;
  wire net_70182_cascademuxed;
  wire net_70188_cascademuxed;
  wire net_7084_cascademuxed;
  wire net_7090_cascademuxed;
  wire net_7096_cascademuxed;
  wire net_7108_cascademuxed;
  wire net_7114_cascademuxed;
  wire net_7120_cascademuxed;
  wire net_7126_cascademuxed;
  wire net_72261_cascademuxed;
  wire net_72267_cascademuxed;
  wire net_72279_cascademuxed;
  wire net_72285_cascademuxed;
  wire net_7231_cascademuxed;
  wire net_7234;
  wire net_72375;
  wire net_72378_cascademuxed;
  wire net_72381;
  wire net_72384_cascademuxed;
  wire net_72387;
  wire net_72390_cascademuxed;
  wire net_72393;
  wire net_72396_cascademuxed;
  wire net_72399;
  wire net_7240;
  wire net_72402_cascademuxed;
  wire net_72405;
  wire net_72408_cascademuxed;
  wire net_72411;
  wire net_72414_cascademuxed;
  wire net_72420_cascademuxed;
  wire net_7246;
  wire net_72501_cascademuxed;
  wire net_7252;
  wire net_72537_cascademuxed;
  wire net_7261_cascademuxed;
  wire net_72624_cascademuxed;
  wire net_72630_cascademuxed;
  wire net_72642_cascademuxed;
  wire net_7273_cascademuxed;
  wire net_72744;
  wire net_72747_cascademuxed;
  wire net_72750;
  wire net_72753_cascademuxed;
  wire net_72756;
  wire net_72759_cascademuxed;
  wire net_72762;
  wire net_72765_cascademuxed;
  wire net_72768;
  wire net_72771_cascademuxed;
  wire net_72774;
  wire net_72777_cascademuxed;
  wire net_72780;
  wire net_72783_cascademuxed;
  wire net_72789_cascademuxed;
  wire net_72870_cascademuxed;
  wire net_72993_cascademuxed;
  wire net_73029_cascademuxed;
  wire net_73113;
  wire net_73116_cascademuxed;
  wire net_73119;
  wire net_73122_cascademuxed;
  wire net_73125;
  wire net_73128_cascademuxed;
  wire net_73131;
  wire net_73134_cascademuxed;
  wire net_73137;
  wire net_73140_cascademuxed;
  wire net_73143;
  wire net_73146_cascademuxed;
  wire net_73275_cascademuxed;
  wire net_73386_cascademuxed;
  wire net_73404_cascademuxed;
  wire net_73497_cascademuxed;
  wire net_73521_cascademuxed;
  wire net_73608_cascademuxed;
  wire net_73626_cascademuxed;
  wire net_73728;
  wire net_73731_cascademuxed;
  wire net_73734;
  wire net_73737_cascademuxed;
  wire net_73740;
  wire net_73743_cascademuxed;
  wire net_73746;
  wire net_73749_cascademuxed;
  wire net_73752;
  wire net_73755_cascademuxed;
  wire net_73758;
  wire net_73761_cascademuxed;
  wire net_73764;
  wire net_73767_cascademuxed;
  wire net_73773_cascademuxed;
  wire net_7384_cascademuxed;
  wire net_73854_cascademuxed;
  wire net_73878_cascademuxed;
  wire net_7390_cascademuxed;
  wire net_7402_cascademuxed;
  wire net_7408_cascademuxed;
  wire net_7543_cascademuxed;
  wire net_7549_cascademuxed;
  wire net_7561_cascademuxed;
  wire net_7861_cascademuxed;
  wire net_79175_cascademuxed;
  wire net_79415_cascademuxed;
  wire net_79538_cascademuxed;
  wire net_79655_cascademuxed;
  wire net_7966_cascademuxed;
  wire net_79679_cascademuxed;
  wire net_79685_cascademuxed;
  wire net_79808_cascademuxed;
  wire net_79937_cascademuxed;
  wire net_80048_cascademuxed;
  wire net_80066_cascademuxed;
  wire net_80177_cascademuxed;
  wire net_80405_cascademuxed;
  wire net_8131_cascademuxed;
  wire net_8143_cascademuxed;
  wire net_8149_cascademuxed;
  wire net_8155_cascademuxed;
  wire net_8266_cascademuxed;
  wire net_83252_cascademuxed;
  wire net_83270_cascademuxed;
  wire net_83399_cascademuxed;
  wire net_83522_cascademuxed;
  wire net_83627_cascademuxed;
  wire net_83729;
  wire net_83732_cascademuxed;
  wire net_83735;
  wire net_83738_cascademuxed;
  wire net_83741;
  wire net_83744_cascademuxed;
  wire net_83747;
  wire net_83750_cascademuxed;
  wire net_83753;
  wire net_83756_cascademuxed;
  wire net_83759;
  wire net_83762_cascademuxed;
  wire net_83765;
  wire net_83768_cascademuxed;
  wire net_83774_cascademuxed;
  wire net_83852;
  wire net_83855_cascademuxed;
  wire net_83858;
  wire net_83861_cascademuxed;
  wire net_83864;
  wire net_83867_cascademuxed;
  wire net_83897_cascademuxed;
  wire net_83990_cascademuxed;
  wire net_8560_cascademuxed;
  wire net_86948_cascademuxed;
  wire net_86960_cascademuxed;
  wire net_86972_cascademuxed;
  wire net_8707_cascademuxed;
  wire net_87083_cascademuxed;
  wire net_87113_cascademuxed;
  wire net_8719_cascademuxed;
  wire net_87218_cascademuxed;
  wire net_87236_cascademuxed;
  wire net_8743_cascademuxed;
  wire net_87563_cascademuxed;
  wire net_87575_cascademuxed;
  wire net_8854_cascademuxed;
  wire net_8866_cascademuxed;
  wire net_9001_cascademuxed;
  wire net_91031_cascademuxed;
  wire net_91067_cascademuxed;
  wire net_9154_cascademuxed;
  wire net_9289_cascademuxed;
  wire net_9295_cascademuxed;
  wire net_9436_cascademuxed;
  wire net_9625_cascademuxed;
  wire net_9748_cascademuxed;
  wire net_9913_cascademuxed;
  wire seg_0_10_sp12_h_r_0_2200;
  wire seg_0_10_sp4_h_r_0_2238;
  wire seg_0_10_sp4_h_r_40_2273;
  wire seg_0_10_sp4_r_v_b_37_2287;
  wire seg_0_10_sp4_r_v_b_39_2289;
  wire seg_0_10_sp4_r_v_b_43_2293;
  wire seg_0_10_sp4_r_v_b_45_2295;
  wire seg_0_10_sp4_r_v_b_47_2297;
  wire seg_0_10_sp4_v_b_11_1454;
  wire seg_0_10_sp4_v_b_16_1656;
  wire seg_0_10_sp4_v_b_18_1658;
  wire seg_0_10_sp4_v_b_3_1446;
  wire seg_0_10_sp4_v_t_36_2298;
  wire seg_0_10_sp4_v_t_47_2309;
  wire seg_0_11_local_g0_1_2315;
  wire seg_0_11_local_g1_0_2322;
  wire seg_0_11_local_g1_5_2327;
  wire seg_0_11_local_g2_0_2330;
  wire seg_0_11_local_g2_1_2331;
  wire seg_0_11_local_g2_2_2332;
  wire seg_0_11_local_g2_3_2333;
  wire seg_0_11_local_g2_4_2334;
  wire seg_0_11_local_g2_6_2336;
  wire seg_0_11_local_g2_7_2337;
  wire seg_0_11_local_g3_0_2338;
  wire seg_0_11_local_g3_1_2339;
  wire seg_0_11_local_g3_2_2340;
  wire seg_0_11_local_g3_4_2342;
  wire seg_0_11_local_g3_5_2343;
  wire seg_0_11_local_g3_7_2345;
  wire seg_0_11_sp12_h_r_1_2407;
  wire seg_0_11_sp4_h_r_0_2444;
  wire seg_0_11_sp4_h_r_10_2446;
  wire seg_0_11_sp4_h_r_12_2448;
  wire seg_0_11_sp4_h_r_13_2449;
  wire seg_0_11_sp4_h_r_17_2453;
  wire seg_0_11_sp4_h_r_26_2463;
  wire seg_0_11_sp4_h_r_2_2456;
  wire seg_0_11_sp4_h_r_30_2468;
  wire seg_0_11_sp4_h_r_31_2469;
  wire seg_0_11_sp4_h_r_33_2471;
  wire seg_0_11_sp4_h_r_34_2472;
  wire seg_0_11_sp4_h_r_35_2473;
  wire seg_0_11_sp4_h_r_46_2485;
  wire seg_0_11_sp4_h_r_47_2486;
  wire seg_0_11_sp4_h_r_4_2478;
  wire seg_0_11_sp4_h_r_6_2488;
  wire seg_0_11_sp4_h_r_7_2489;
  wire seg_0_11_sp4_h_r_8_2490;
  wire seg_0_11_sp4_h_r_9_2491;
  wire seg_0_11_sp4_r_v_b_0_1850;
  wire seg_0_11_sp4_r_v_b_12_2076;
  wire seg_0_11_sp4_r_v_b_16_2080;
  wire seg_0_11_sp4_r_v_b_20_2084;
  wire seg_0_11_sp4_r_v_b_8_1858;
  wire seg_0_11_sp4_v_b_29_2092;
  wire seg_0_11_sp4_v_b_33_2096;
  wire seg_0_11_sp4_v_b_4_1657;
  wire seg_0_11_sp4_v_b_5_1656;
  wire seg_0_11_sp4_v_b_7_1658;
  wire seg_0_12_local_g0_0_2520;
  wire seg_0_12_local_g0_1_2521;
  wire seg_0_12_local_g0_2_2522;
  wire seg_0_12_local_g0_3_2523;
  wire seg_0_12_local_g0_4_2524;
  wire seg_0_12_local_g0_6_2526;
  wire seg_0_12_local_g1_0_2528;
  wire seg_0_12_local_g1_1_2529;
  wire seg_0_12_local_g1_2_2530;
  wire seg_0_12_local_g1_3_2531;
  wire seg_0_12_local_g1_5_2533;
  wire seg_0_12_local_g1_6_2534;
  wire seg_0_12_local_g1_7_2535;
  wire seg_0_12_local_g3_0_2544;
  wire seg_0_12_local_g3_2_2546;
  wire seg_0_12_local_g3_4_2548;
  wire seg_0_12_sp12_h_r_0_2614;
  wire seg_0_12_sp12_h_r_6_2634;
  wire seg_0_12_sp4_h_r_10_2654;
  wire seg_0_12_sp4_h_r_11_2655;
  wire seg_0_12_sp4_h_r_16_2660;
  wire seg_0_12_sp4_h_r_20_2665;
  wire seg_0_12_sp4_h_r_28_2673;
  wire seg_0_12_sp4_h_r_2_2664;
  wire seg_0_12_sp4_h_r_4_2686;
  wire seg_0_12_sp4_r_v_b_11_2086;
  wire seg_0_12_sp4_r_v_b_25_2492;
  wire seg_0_12_sp4_r_v_b_31_2498;
  wire seg_0_12_sp4_r_v_b_39_2703;
  wire seg_0_12_sp4_v_b_12_2088;
  wire seg_0_12_sp4_v_b_13_2089;
  wire seg_0_12_sp4_v_b_17_2093;
  wire seg_0_12_sp4_v_b_19_2095;
  wire seg_0_12_sp4_v_b_1_1861;
  wire seg_0_12_sp4_v_b_24_2299;
  wire seg_0_12_sp4_v_b_34_2309;
  wire seg_0_12_sp4_v_b_42_2510;
  wire seg_0_12_sp4_v_b_4_1866;
  wire seg_0_12_sp4_v_b_6_1868;
  wire seg_0_12_sp4_v_b_7_1867;
  wire seg_0_12_sp4_v_b_8_1870;
  wire seg_0_12_sp4_v_t_43_2719;
  wire seg_0_12_sp4_v_t_45_2721;
  wire seg_0_13_sp4_h_r_0_2861;
  wire seg_0_13_sp4_h_r_24_2878;
  wire seg_0_13_sp4_h_r_38_2893;
  wire seg_0_13_sp4_h_r_4_2895;
  wire seg_0_13_sp4_h_r_8_2907;
  wire seg_0_13_sp4_r_v_b_21_2501;
  wire seg_0_13_sp4_r_v_b_27_2702;
  wire seg_0_13_sp4_r_v_b_3_2288;
  wire seg_0_13_sp4_v_b_11_2098;
  wire seg_0_13_sp4_v_b_12_2298;
  wire seg_0_13_sp4_v_b_2_2091;
  wire seg_0_13_sp4_v_b_3_2090;
  wire seg_0_13_sp4_v_b_7_2094;
  wire seg_0_13_sp4_v_b_8_2097;
  wire seg_0_14_sp4_v_b_11_2308;
  wire seg_0_14_sp4_v_b_7_2304;
  wire seg_0_14_sp4_v_t_39_3151;
  wire seg_0_14_sp4_v_t_45_3157;
  wire seg_0_14_sp4_v_t_46_3158;
  wire seg_0_15_sp4_h_r_10_3300;
  wire seg_0_15_sp4_h_r_14_3304;
  wire seg_0_15_sp4_h_r_16_3306;
  wire seg_0_15_sp4_h_r_18_3308;
  wire seg_0_15_sp4_h_r_8_3344;
  wire seg_0_15_sp4_r_v_b_23_2920;
  wire seg_0_15_sp4_v_b_20_2720;
  wire seg_0_15_sp4_v_b_28_2926;
  wire seg_0_15_sp4_v_t_40_3362;
  wire seg_0_15_sp4_v_t_43_3365;
  wire seg_0_16_local_g0_6_3380;
  wire seg_0_16_local_g1_0_3382;
  wire seg_0_16_local_g1_1_3383;
  wire seg_0_16_local_g1_3_3385;
  wire seg_0_16_local_g1_4_3386;
  wire seg_0_16_local_g1_6_3388;
  wire seg_0_16_local_g1_7_3389;
  wire seg_0_16_local_g2_0_3390;
  wire seg_0_16_local_g2_2_3392;
  wire seg_0_16_local_g2_3_3393;
  wire seg_0_16_local_g2_4_3394;
  wire seg_0_16_local_g2_5_3395;
  wire seg_0_16_local_g2_7_3397;
  wire seg_0_16_local_g3_1_3399;
  wire seg_0_16_local_g3_2_3400;
  wire seg_0_16_local_g3_4_3402;
  wire seg_0_16_sp12_v_b_10_2014;
  wire seg_0_16_sp4_h_r_18_3514;
  wire seg_0_16_sp4_h_r_28_3525;
  wire seg_0_16_sp4_h_r_31_3529;
  wire seg_0_16_sp4_h_r_33_3531;
  wire seg_0_16_sp4_h_r_45_3544;
  wire seg_0_16_sp4_r_v_b_0_2910;
  wire seg_0_16_sp4_r_v_b_11_2919;
  wire seg_0_16_sp4_r_v_b_13_3137;
  wire seg_0_16_sp4_r_v_b_15_3139;
  wire seg_0_16_sp4_r_v_b_18_3142;
  wire seg_0_16_sp4_r_v_b_1_2909;
  wire seg_0_16_sp4_r_v_b_3_2911;
  wire seg_0_16_sp4_r_v_b_44_3560;
  wire seg_0_16_sp4_r_v_b_4_2914;
  wire seg_0_16_sp4_r_v_b_5_2913;
  wire seg_0_16_sp4_r_v_b_6_2916;
  wire seg_0_16_sp4_r_v_b_8_2918;
  wire seg_0_16_sp4_v_b_10_2723;
  wire seg_0_16_sp4_v_b_22_2931;
  wire seg_0_16_sp4_v_b_23_2932;
  wire seg_0_16_sp4_v_b_26_3151;
  wire seg_0_16_sp4_v_b_32_3157;
  wire seg_0_16_sp4_v_b_6_2719;
  wire seg_0_16_sp4_v_b_8_2721;
  wire seg_0_16_sp4_v_b_9_2720;
  wire seg_0_17_local_g0_0_3580;
  wire seg_0_17_local_g0_2_3582;
  wire seg_0_17_local_g0_3_3583;
  wire seg_0_17_local_g0_5_3585;
  wire seg_0_17_local_g0_7_3587;
  wire seg_0_17_local_g1_1_3589;
  wire seg_0_17_local_g1_2_3590;
  wire seg_0_17_local_g1_4_3592;
  wire seg_0_17_local_g1_6_3594;
  wire seg_0_17_local_g1_7_3595;
  wire seg_0_17_local_g2_1_3597;
  wire seg_0_17_local_g2_2_3598;
  wire seg_0_17_local_g2_4_3600;
  wire seg_0_17_local_g3_2_3606;
  wire seg_0_17_local_g3_3_3607;
  wire seg_0_17_local_g3_7_3611;
  wire seg_0_17_sp4_h_r_0_3712;
  wire seg_0_17_sp4_h_r_18_3722;
  wire seg_0_17_sp4_h_r_26_3731;
  wire seg_0_17_sp4_h_r_2_3724;
  wire seg_0_17_sp4_h_r_4_3746;
  wire seg_0_17_sp4_h_r_6_3756;
  wire seg_0_17_sp4_h_r_8_3758;
  wire seg_0_17_sp4_r_v_b_10_3147;
  wire seg_0_17_sp4_r_v_b_12_3346;
  wire seg_0_17_sp4_r_v_b_17_3351;
  wire seg_0_17_sp4_r_v_b_18_3352;
  wire seg_0_17_sp4_r_v_b_19_3353;
  wire seg_0_17_sp4_r_v_b_1_3136;
  wire seg_0_17_sp4_r_v_b_23_3357;
  wire seg_0_17_sp4_r_v_b_28_3557;
  wire seg_0_17_sp4_r_v_b_29_3556;
  wire seg_0_17_sp4_r_v_b_31_3558;
  wire seg_0_17_sp4_r_v_b_35_3562;
  wire seg_0_17_sp4_r_v_b_9_3144;
  wire seg_0_17_sp4_v_b_18_3154;
  wire seg_0_17_sp4_v_b_22_3158;
  wire seg_0_17_sp4_v_b_23_3159;
  wire seg_0_17_sp4_v_b_2_2924;
  wire seg_0_17_sp4_v_b_30_3365;
  wire seg_0_17_sp4_v_b_3_2923;
  wire seg_0_17_sp4_v_b_4_2926;
  wire seg_0_17_sp4_v_b_5_2925;
  wire seg_0_17_sp4_v_b_6_2928;
  wire seg_0_17_sp4_v_b_8_2930;
  wire seg_0_18_sp4_h_r_6_3965;
  wire seg_0_18_sp4_r_v_b_11_3356;
  wire seg_0_18_sp4_r_v_b_13_3553;
  wire seg_0_18_sp4_r_v_b_19_3559;
  wire seg_0_18_sp4_r_v_b_5_3350;
  wire seg_0_18_sp4_r_v_b_9_3354;
  wire seg_0_18_sp4_v_b_16_3362;
  wire seg_0_19_sp12_v_b_1_1578;
  wire seg_0_20_sp12_v_b_1_1787;
  wire seg_0_20_sp4_v_b_10_3575;
  wire seg_0_20_sp4_v_t_36_4435;
  wire seg_0_21_sp12_v_b_5_2430;
  wire seg_0_21_sp4_h_r_0_4602;
  wire seg_0_21_sp4_h_r_1_4603;
  wire seg_0_21_sp4_h_r_2_4614;
  wire seg_0_21_sp4_h_r_4_4636;
  wire seg_0_21_sp4_v_b_0_3773;
  wire seg_0_21_sp4_v_b_1_3772;
  wire seg_0_21_sp4_v_b_2_3775;
  wire seg_0_21_sp4_v_b_5_3776;
  wire seg_0_21_sp4_v_b_6_3779;
  wire seg_0_22_sp12_v_b_0_2225;
  wire seg_0_22_sp4_h_r_0_4829;
  wire seg_0_22_sp4_h_r_8_4875;
  wire seg_0_22_sp4_v_b_3_3983;
  wire seg_0_22_sp4_v_t_47_4900;
  wire seg_0_23_sp4_h_r_0_5039;
  wire seg_0_23_sp4_r_v_b_11_4433;
  wire seg_0_23_sp4_r_v_b_15_4653;
  wire seg_0_23_sp4_r_v_b_3_4425;
  wire seg_0_23_sp4_r_v_b_5_4427;
  wire seg_0_23_sp4_r_v_b_7_4429;
  wire seg_0_23_sp4_r_v_b_9_4431;
  wire seg_0_23_sp4_v_b_12_4435;
  wire seg_0_24_local_g0_2_5117;
  wire seg_0_24_local_g0_3_5118;
  wire seg_0_24_local_g0_5_5120;
  wire seg_0_24_local_g0_7_5122;
  wire seg_0_24_local_g1_0_5123;
  wire seg_0_24_local_g1_2_5125;
  wire seg_0_24_local_g1_3_5126;
  wire seg_0_24_local_g1_4_5127;
  wire seg_0_24_local_g1_5_5128;
  wire seg_0_24_local_g2_2_5133;
  wire seg_0_24_local_g2_3_5134;
  wire seg_0_24_local_g3_1_5140;
  wire seg_0_24_local_g3_2_5141;
  wire seg_0_24_local_g3_3_5142;
  wire seg_0_24_local_g3_5_5144;
  wire seg_0_24_local_g3_7_5146;
  wire seg_0_24_sp4_h_r_12_5249;
  wire seg_0_24_sp4_h_r_18_5255;
  wire seg_0_24_sp4_h_r_22_5260;
  wire seg_0_24_sp4_h_r_35_5274;
  wire seg_0_24_sp4_r_v_b_11_4660;
  wire seg_0_24_sp4_r_v_b_15_4880;
  wire seg_0_24_sp4_r_v_b_17_4882;
  wire seg_0_24_sp4_r_v_b_18_4883;
  wire seg_0_24_sp4_r_v_b_19_4884;
  wire seg_0_24_sp4_r_v_b_1_4650;
  wire seg_0_24_sp4_r_v_b_21_4886;
  wire seg_0_24_sp4_r_v_b_23_4888;
  wire seg_0_24_sp4_r_v_b_27_5089;
  wire seg_0_24_sp4_r_v_b_29_5091;
  wire seg_0_24_sp4_r_v_b_34_5098;
  wire seg_0_24_sp4_r_v_b_35_5097;
  wire seg_0_24_sp4_r_v_b_5_4654;
  wire seg_0_24_sp4_r_v_b_9_4658;
  wire seg_0_24_sp4_v_b_10_4446;
  wire seg_0_24_sp4_v_b_13_4663;
  wire seg_0_24_sp4_v_b_16_4666;
  wire seg_0_24_sp4_v_b_19_4669;
  wire seg_0_24_sp4_v_b_21_4671;
  wire seg_0_24_sp4_v_b_23_4673;
  wire seg_0_25_local_g0_2_5323;
  wire seg_0_25_local_g0_4_5325;
  wire seg_0_25_local_g0_5_5326;
  wire seg_0_25_local_g0_6_5327;
  wire seg_0_25_local_g0_7_5328;
  wire seg_0_25_local_g1_0_5329;
  wire seg_0_25_local_g1_1_5330;
  wire seg_0_25_local_g1_2_5331;
  wire seg_0_25_local_g1_3_5332;
  wire seg_0_25_local_g1_7_5336;
  wire seg_0_25_local_g2_3_5340;
  wire seg_0_25_local_g2_4_5341;
  wire seg_0_25_local_g2_5_5342;
  wire seg_0_25_local_g2_7_5344;
  wire seg_0_25_local_g3_0_5345;
  wire seg_0_25_local_g3_1_5346;
  wire seg_0_25_sp12_h_r_2_5427;
  wire seg_0_25_sp12_h_r_3_5432;
  wire seg_0_25_sp12_v_b_13_4134;
  wire seg_0_25_sp12_v_b_19_4816;
  wire seg_0_25_sp4_h_r_0_5453;
  wire seg_0_25_sp4_h_r_24_5470;
  wire seg_0_25_sp4_h_r_26_5472;
  wire seg_0_25_sp4_h_r_6_5497;
  wire seg_0_25_sp4_h_r_8_5499;
  wire seg_0_25_sp4_r_v_b_0_4878;
  wire seg_0_25_sp4_r_v_b_12_5087;
  wire seg_0_25_sp4_r_v_b_13_5088;
  wire seg_0_25_sp4_r_v_b_15_5090;
  wire seg_0_25_sp4_r_v_b_17_5092;
  wire seg_0_25_sp4_r_v_b_31_5299;
  wire seg_0_25_sp4_r_v_b_3_4879;
  wire seg_0_25_sp4_r_v_b_5_4881;
  wire seg_0_25_sp4_v_b_13_4890;
  wire seg_0_25_sp4_v_b_14_4891;
  wire seg_0_25_sp4_v_b_15_4892;
  wire seg_0_25_sp4_v_b_2_4665;
  wire seg_0_25_sp4_v_b_4_4667;
  wire seg_0_25_sp4_v_b_7_4668;
  wire seg_0_25_sp4_v_b_9_4670;
  wire seg_0_26_sp4_h_r_28_5683;
  wire seg_0_26_sp4_r_v_b_17_5298;
  wire seg_0_26_sp4_r_v_b_21_5302;
  wire seg_0_26_sp4_r_v_b_35_5511;
  wire seg_0_26_sp4_r_v_b_7_5093;
  wire seg_0_26_sp4_r_v_b_9_5095;
  wire seg_0_26_sp4_v_b_10_4900;
  wire seg_0_4_sp4_v_t_39_1031;
  wire seg_0_4_sp4_v_t_45_1037;
  wire seg_0_5_sp4_h_r_0_1178;
  wire seg_0_5_sp4_h_r_11_1181;
  wire seg_0_5_sp4_h_r_14_1184;
  wire seg_0_5_sp4_h_r_24_1195;
  wire seg_0_5_sp4_h_r_28_1199;
  wire seg_0_5_sp4_h_r_34_1206;
  wire seg_0_5_sp4_h_r_38_1210;
  wire seg_0_5_sp4_h_r_3_1201;
  wire seg_0_5_sp4_h_r_7_1223;
  wire seg_0_5_sp4_h_r_8_1224;
  wire seg_0_5_sp4_r_v_b_21_798;
  wire seg_0_5_sp4_v_b_26_804;
  wire seg_0_5_sp4_v_t_36_1238;
  wire seg_0_6_local_g0_3_1257;
  wire seg_0_6_local_g0_4_1258;
  wire seg_0_6_local_g0_5_1259;
  wire seg_0_6_local_g1_0_1262;
  wire seg_0_6_local_g1_2_1264;
  wire seg_0_6_local_g1_5_1267;
  wire seg_0_6_local_g1_6_1268;
  wire seg_0_6_local_g2_2_1272;
  wire seg_0_6_local_g2_4_1274;
  wire seg_0_6_local_g2_5_1275;
  wire seg_0_6_local_g2_6_1276;
  wire seg_0_6_local_g3_0_1278;
  wire seg_0_6_local_g3_1_1279;
  wire seg_0_6_local_g3_2_1280;
  wire seg_0_6_local_g3_3_1281;
  wire seg_0_6_local_g3_7_1285;
  wire seg_0_6_sp4_h_r_0_1384;
  wire seg_0_6_sp4_h_r_29_1406;
  wire seg_0_6_sp4_h_r_42_1421;
  wire seg_0_6_sp4_h_r_44_1423;
  wire seg_0_6_sp4_h_r_4_1418;
  wire seg_0_6_sp4_h_r_5_1427;
  wire seg_0_6_sp4_h_r_8_1430;
  wire seg_0_6_sp4_h_r_9_1431;
  wire seg_0_6_sp4_r_v_b_14_1018;
  wire seg_0_6_sp4_r_v_b_15_1019;
  wire seg_0_6_sp4_r_v_b_16_1020;
  wire seg_0_6_sp4_r_v_b_19_1023;
  wire seg_0_6_sp4_r_v_b_27_1228;
  wire seg_0_6_sp4_r_v_b_36_1432;
  wire seg_0_6_sp4_r_v_b_41_1437;
  wire seg_0_6_sp4_r_v_b_42_1438;
  wire seg_0_6_sp4_r_v_b_43_1439;
  wire seg_0_6_sp4_v_b_12_801;
  wire seg_0_6_sp4_v_b_13_802;
  wire seg_0_6_sp4_v_b_14_803;
  wire seg_0_6_sp4_v_b_16_805;
  wire seg_0_6_sp4_v_b_18_807;
  wire seg_0_6_sp4_v_b_19_808;
  wire seg_0_6_sp4_v_b_21_810;
  wire seg_0_6_sp4_v_b_22_811;
  wire seg_0_6_sp4_v_b_39_1241;
  wire seg_0_6_sp4_v_t_39_1447;
  wire seg_0_7_local_g0_1_1461;
  wire seg_0_7_local_g0_4_1464;
  wire seg_0_7_local_g1_3_1471;
  wire seg_0_7_local_g1_6_1474;
  wire seg_0_7_local_g2_0_1476;
  wire seg_0_7_local_g2_2_1478;
  wire seg_0_7_local_g2_3_1479;
  wire seg_0_7_local_g2_7_1483;
  wire seg_0_7_local_g3_0_1484;
  wire seg_0_7_local_g3_1_1485;
  wire seg_0_7_local_g3_2_1486;
  wire seg_0_7_local_g3_3_1487;
  wire seg_0_7_local_g3_4_1488;
  wire seg_0_7_local_g3_5_1489;
  wire seg_0_7_local_g3_6_1490;
  wire seg_0_7_local_g3_7_1491;
  wire seg_0_7_neigh_op_bnr_3_1133;
  wire seg_0_7_neigh_op_bnr_6_1136;
  wire seg_0_7_neigh_op_tnr_3_1547;
  wire seg_0_7_neigh_op_tnr_4_1548;
  wire seg_0_7_neigh_op_tnr_7_1551;
  wire seg_0_7_sp12_h_r_1_1555;
  wire seg_0_7_sp4_h_r_0_1592;
  wire seg_0_7_sp4_h_r_10_1594;
  wire seg_0_7_sp4_h_r_12_1596;
  wire seg_0_7_sp4_h_r_14_1598;
  wire seg_0_7_sp4_h_r_17_1601;
  wire seg_0_7_sp4_h_r_1_1593;
  wire seg_0_7_sp4_h_r_25_1610;
  wire seg_0_7_sp4_h_r_32_1618;
  wire seg_0_7_sp4_h_r_3_1615;
  wire seg_0_7_sp4_h_r_40_1627;
  wire seg_0_7_sp4_h_r_47_1634;
  wire seg_0_7_sp4_h_r_4_1626;
  wire seg_0_7_sp4_h_r_6_1636;
  wire seg_0_7_sp4_h_r_7_1637;
  wire seg_0_7_sp4_h_r_8_1638;
  wire seg_0_7_sp4_r_v_b_13_1227;
  wire seg_0_7_sp4_r_v_b_19_1233;
  wire seg_0_7_sp4_r_v_b_21_1235;
  wire seg_0_7_sp4_r_v_b_22_1236;
  wire seg_0_7_sp4_r_v_b_34_1443;
  wire seg_0_7_sp4_r_v_b_41_1645;
  wire seg_0_7_sp4_r_v_b_42_1646;
  wire seg_0_7_sp4_r_v_b_45_1649;
  wire seg_0_7_sp4_v_b_11_811;
  wire seg_0_7_sp4_v_b_2_804;
  wire seg_0_7_sp4_v_b_35_1248;
  wire seg_0_7_sp4_v_b_40_1448;
  wire seg_0_7_sp4_v_t_37_1653;
  wire seg_0_7_sp4_v_t_44_1660;
  wire seg_0_8_sp12_h_r_1_1764;
  wire seg_0_8_sp4_h_r_0_1801;
  wire seg_0_8_sp4_h_r_10_1803;
  wire seg_0_8_sp4_h_r_12_1805;
  wire seg_0_8_sp4_h_r_1_1802;
  wire seg_0_8_sp4_h_r_20_1814;
  wire seg_0_8_sp4_h_r_2_1813;
  wire seg_0_8_sp4_h_r_6_1845;
  wire seg_0_8_sp4_h_r_7_1846;
  wire seg_0_8_sp4_r_v_b_7_1232;
  wire seg_0_8_sp4_v_b_26_1447;
  wire seg_0_8_sp4_v_b_2_1031;
  wire seg_0_8_sp4_v_b_8_1037;
  wire seg_0_9_sp12_h_r_1_1991;
  wire seg_0_9_sp4_h_r_0_2028;
  wire seg_0_9_sp4_h_r_10_2030;
  wire seg_0_9_sp4_h_r_11_2031;
  wire seg_0_9_sp4_h_r_2_2040;
  wire seg_0_9_sp4_h_r_5_2071;
  wire seg_0_9_sp4_h_r_6_2072;
  wire seg_0_9_sp4_h_r_9_2075;
  wire seg_0_9_sp4_v_b_11_1248;
  wire seg_0_9_sp4_v_b_3_1240;
  wire seg_0_9_sp4_v_b_7_1244;
  wire seg_0_9_sp4_v_b_8_1247;
  wire seg_0_9_sp4_v_t_36_2088;
  wire seg_10_10_glb_netwk_0_5;
  wire seg_10_10_glb_netwk_4_9;
  wire seg_10_10_local_g0_1_42436;
  wire seg_10_10_local_g0_2_42437;
  wire seg_10_10_local_g0_4_42439;
  wire seg_10_10_local_g1_1_42444;
  wire seg_10_10_local_g1_2_42445;
  wire seg_10_10_local_g1_5_42448;
  wire seg_10_10_local_g2_3_42454;
  wire seg_10_10_local_g2_5_42456;
  wire seg_10_10_lutff_1_out_38564;
  wire seg_10_10_lutff_3_out_38566;
  wire seg_10_10_lutff_5_out_38568;
  wire seg_10_10_sp12_h_r_1_42526;
  wire seg_10_10_sp12_h_r_20_2200;
  wire seg_10_10_sp4_h_l_39_27629;
  wire seg_10_10_sp4_h_l_41_27631;
  wire seg_10_10_sp4_h_l_43_27633;
  wire seg_10_10_sp4_h_r_0_42529;
  wire seg_10_10_sp4_h_r_14_38703;
  wire seg_10_10_sp4_h_r_18_38707;
  wire seg_10_10_sp4_h_r_28_34873;
  wire seg_10_10_sp4_h_r_32_34877;
  wire seg_10_10_sp4_h_r_3_42534;
  wire seg_10_10_sp4_h_r_4_42535;
  wire seg_10_10_sp4_r_v_b_29_42422;
  wire seg_10_10_sp4_v_b_14_38466;
  wire seg_10_10_sp4_v_b_20_38472;
  wire seg_10_10_sp4_v_b_2_38344;
  wire seg_10_10_sp4_v_b_32_38596;
  wire seg_10_10_sp4_v_b_46_38720;
  wire seg_10_10_sp4_v_b_4_38346;
  wire seg_10_10_sp4_v_t_46_38843;
  wire seg_10_11_glb_netwk_0_5;
  wire seg_10_11_local_g0_0_42558;
  wire seg_10_11_local_g0_1_42559;
  wire seg_10_11_local_g0_2_42560;
  wire seg_10_11_local_g0_7_42565;
  wire seg_10_11_local_g1_1_42567;
  wire seg_10_11_local_g1_3_42569;
  wire seg_10_11_local_g1_6_42572;
  wire seg_10_11_local_g2_1_42575;
  wire seg_10_11_local_g2_2_42576;
  wire seg_10_11_local_g2_7_42581;
  wire seg_10_11_local_g3_6_42588;
  wire seg_10_11_lutff_0_out_38686;
  wire seg_10_11_lutff_1_out_38687;
  wire seg_10_11_lutff_3_out_38689;
  wire seg_10_11_lutff_6_out_38692;
  wire seg_10_11_neigh_op_bnr_1_42395;
  wire seg_10_11_neigh_op_bnr_7_42401;
  wire seg_10_11_sp4_h_r_17_38827;
  wire seg_10_11_sp4_h_r_1_42653;
  wire seg_10_11_sp4_h_r_24_34990;
  wire seg_10_11_sp4_h_r_26_34994;
  wire seg_10_11_sp4_h_r_30_34998;
  wire seg_10_11_sp4_h_r_31_34999;
  wire seg_10_11_sp4_r_v_b_22_42428;
  wire seg_10_11_sp4_r_v_b_26_42544;
  wire seg_10_11_sp4_r_v_b_33_42549;
  wire seg_10_11_sp4_r_v_b_6_42302;
  wire seg_10_11_sp4_v_b_3_38466;
  wire seg_10_11_sp4_v_b_5_38468;
  wire seg_10_12_glb_netwk_0_5;
  wire seg_10_12_local_g0_2_42683;
  wire seg_10_12_local_g1_3_42692;
  wire seg_10_12_sp12_v_b_0_41270;
  wire seg_10_12_sp4_h_r_11_42778;
  wire seg_10_12_sp4_h_r_20_38955;
  wire seg_10_12_sp4_v_b_0_38588;
  wire seg_10_12_sp4_v_b_18_38716;
  wire seg_10_12_sp4_v_b_1_38587;
  wire seg_10_12_sp4_v_b_3_38589;
  wire seg_10_12_sp4_v_b_6_38594;
  wire seg_10_12_sp4_v_b_7_38593;
  wire seg_10_12_sp4_v_b_8_38596;
  wire seg_10_13_glb_netwk_0_5;
  wire seg_10_13_local_g0_2_42806;
  wire seg_10_13_local_g0_6_42810;
  wire seg_10_13_local_g1_2_42814;
  wire seg_10_13_lutff_1_out_38933;
  wire seg_10_13_lutff_2_out_38934;
  wire seg_10_13_sp4_h_l_36_27932;
  wire seg_10_13_sp4_h_r_14_39072;
  wire seg_10_13_sp4_h_r_9_42909;
  wire seg_10_13_sp4_r_v_b_26_42790;
  wire seg_10_13_sp4_v_b_0_38711;
  wire seg_10_13_sp4_v_b_1_38710;
  wire seg_10_13_sp4_v_b_2_38713;
  wire seg_10_13_sp4_v_b_9_38718;
  wire seg_10_13_sp4_v_t_46_39212;
  wire seg_10_14_glb_netwk_0_5;
  wire seg_10_14_local_g0_0_42927;
  wire seg_10_14_local_g1_1_42936;
  wire seg_10_14_local_g3_0_42951;
  wire seg_10_14_local_g3_1_42952;
  wire seg_10_14_local_g3_2_42953;
  wire seg_10_14_local_g3_3_42954;
  wire seg_10_14_local_g3_4_42955;
  wire seg_10_14_sp4_h_l_46_28036;
  wire seg_10_14_sp4_h_r_10_43023;
  wire seg_10_14_sp4_h_r_16_39197;
  wire seg_10_14_sp4_h_r_24_35359;
  wire seg_10_14_sp4_h_r_35_35362;
  wire seg_10_14_sp4_h_r_3_43026;
  wire seg_10_14_sp4_r_v_b_17_42792;
  wire seg_10_14_sp4_r_v_b_19_42794;
  wire seg_10_14_sp4_r_v_b_20_42795;
  wire seg_10_14_sp4_r_v_b_23_42798;
  wire seg_10_14_sp4_r_v_b_40_43037;
  wire seg_10_14_sp4_r_v_b_42_43039;
  wire seg_10_14_sp4_v_b_14_38958;
  wire seg_10_14_sp4_v_b_16_38960;
  wire seg_10_14_sp4_v_b_9_38841;
  wire seg_10_15_glb_netwk_0_5;
  wire seg_10_15_local_g0_2_43052;
  wire seg_10_15_local_g0_3_43053;
  wire seg_10_15_local_g0_6_43056;
  wire seg_10_15_local_g1_3_43061;
  wire seg_10_15_local_g1_5_43063;
  wire seg_10_15_local_g1_7_43065;
  wire seg_10_15_local_g3_2_43076;
  wire seg_10_15_local_g3_3_43077;
  wire seg_10_15_lutff_0_out_39178;
  wire seg_10_15_lutff_4_out_39182;
  wire seg_10_15_lutff_7_out_39185;
  wire seg_10_15_neigh_op_bnl_2_35226;
  wire seg_10_15_sp4_h_l_36_28136;
  wire seg_10_15_sp4_h_l_43_28143;
  wire seg_10_15_sp4_h_r_10_43146;
  wire seg_10_15_sp4_h_r_18_39322;
  wire seg_10_15_sp4_h_r_2_43148;
  wire seg_10_15_sp4_r_v_b_27_43035;
  wire seg_10_15_sp4_r_v_b_29_43037;
  wire seg_10_15_sp4_v_b_11_38966;
  wire seg_10_15_sp4_v_b_22_39089;
  wire seg_10_15_sp4_v_b_35_39212;
  wire seg_10_15_sp4_v_b_36_39325;
  wire seg_10_15_sp4_v_b_3_38958;
  wire seg_10_16_glb_netwk_0_5;
  wire seg_10_16_local_g1_1_43182;
  wire seg_10_16_local_g1_6_43187;
  wire seg_10_16_local_g2_2_43191;
  wire seg_10_16_local_g2_3_43192;
  wire seg_10_16_local_g2_4_43193;
  wire seg_10_16_local_g2_7_43196;
  wire seg_10_16_lutff_0_out_39301;
  wire seg_10_16_lutff_1_out_39302;
  wire seg_10_16_lutff_3_out_39304;
  wire seg_10_16_lutff_4_out_39305;
  wire seg_10_16_lutff_5_out_39306;
  wire seg_10_16_sp12_h_r_9_28234;
  wire seg_10_16_sp12_v_b_7_42159;
  wire seg_10_16_sp4_h_r_22_39439;
  wire seg_10_16_sp4_h_r_26_35609;
  wire seg_10_16_sp4_h_r_3_43272;
  wire seg_10_16_sp4_h_r_7_43276;
  wire seg_10_16_sp4_r_v_b_12_43033;
  wire seg_10_16_sp4_v_b_27_39327;
  wire seg_10_16_sp4_v_b_2_39082;
  wire seg_10_16_sp4_v_b_8_39088;
  wire seg_10_16_sp4_v_t_46_39581;
  wire seg_10_17_glb_netwk_0_5;
  wire seg_10_17_local_g0_0_43296;
  wire seg_10_17_local_g0_2_43298;
  wire seg_10_17_local_g0_3_43299;
  wire seg_10_17_local_g0_4_43300;
  wire seg_10_17_local_g0_5_43301;
  wire seg_10_17_local_g0_6_43302;
  wire seg_10_17_local_g1_1_43305;
  wire seg_10_17_local_g1_3_43307;
  wire seg_10_17_local_g1_6_43310;
  wire seg_10_17_local_g2_3_43315;
  wire seg_10_17_local_g2_4_43316;
  wire seg_10_17_local_g2_7_43319;
  wire seg_10_17_lutff_0_out_39424;
  wire seg_10_17_lutff_1_out_39425;
  wire seg_10_17_lutff_2_out_39426;
  wire seg_10_17_lutff_4_out_39428;
  wire seg_10_17_lutff_6_out_39430;
  wire seg_10_17_lutff_7_out_39431;
  wire seg_10_17_neigh_op_bot_0_39301;
  wire seg_10_17_neigh_op_bot_4_39305;
  wire seg_10_17_neigh_op_bot_5_39306;
  wire seg_10_17_neigh_op_rgt_3_43258;
  wire seg_10_17_neigh_op_rgt_4_43259;
  wire seg_10_17_neigh_op_rgt_7_43262;
  wire seg_10_17_sp4_h_r_11_43393;
  wire seg_10_17_sp4_h_r_18_39568;
  wire seg_10_17_sp4_h_r_22_39562;
  wire seg_10_17_sp4_r_v_b_1_43033;
  wire seg_10_17_sp4_r_v_b_3_43035;
  wire seg_10_17_sp4_v_b_0_39203;
  wire seg_10_17_sp4_v_b_14_39327;
  wire seg_10_17_sp4_v_b_4_39207;
  wire seg_10_18_glb_netwk_0_5;
  wire seg_10_18_glb_netwk_1_6;
  wire seg_10_18_glb_netwk_4_9;
  wire seg_10_18_local_g0_0_43419;
  wire seg_10_18_local_g0_2_43421;
  wire seg_10_18_local_g0_3_43422;
  wire seg_10_18_local_g0_6_43425;
  wire seg_10_18_local_g0_7_43426;
  wire seg_10_18_local_g1_1_43428;
  wire seg_10_18_local_g1_4_43431;
  wire seg_10_18_local_g1_5_43432;
  wire seg_10_18_local_g1_7_43434;
  wire seg_10_18_local_g2_0_43435;
  wire seg_10_18_local_g2_2_43437;
  wire seg_10_18_local_g2_3_43438;
  wire seg_10_18_local_g2_4_43439;
  wire seg_10_18_local_g2_6_43441;
  wire seg_10_18_local_g3_1_43444;
  wire seg_10_18_local_g3_5_43448;
  wire seg_10_18_local_g3_7_43450;
  wire seg_10_18_lutff_1_out_39548;
  wire seg_10_18_lutff_2_out_39549;
  wire seg_10_18_lutff_3_out_39550;
  wire seg_10_18_lutff_5_out_39552;
  wire seg_10_18_lutff_6_out_39553;
  wire seg_10_18_lutff_7_out_39554;
  wire seg_10_18_neigh_op_lft_0_35716;
  wire seg_10_18_neigh_op_lft_2_35718;
  wire seg_10_18_neigh_op_lft_5_35721;
  wire seg_10_18_neigh_op_lft_6_35722;
  wire seg_10_18_neigh_op_lft_7_35723;
  wire seg_10_18_neigh_op_rgt_1_43379;
  wire seg_10_18_sp4_h_r_0_43513;
  wire seg_10_18_sp4_h_r_3_43518;
  wire seg_10_18_sp4_h_r_8_43523;
  wire seg_10_18_sp4_r_v_b_12_43279;
  wire seg_10_18_sp4_r_v_b_4_43161;
  wire seg_10_18_sp4_r_v_b_8_43165;
  wire seg_10_18_sp4_v_b_31_39577;
  wire seg_10_19_glb_netwk_0_5;
  wire seg_10_19_glb_netwk_4_9;
  wire seg_10_19_local_g0_2_43544;
  wire seg_10_19_local_g0_7_43549;
  wire seg_10_19_local_g1_1_43551;
  wire seg_10_19_local_g1_6_43556;
  wire seg_10_19_local_g1_7_43557;
  wire seg_10_19_local_g2_1_43559;
  wire seg_10_19_local_g3_2_43568;
  wire seg_10_19_local_g3_3_43569;
  wire seg_10_19_neigh_op_rgt_1_43502;
  wire seg_10_19_sp12_v_b_11_42774;
  wire seg_10_19_sp12_v_b_2_42281;
  wire seg_10_19_sp4_h_r_18_39814;
  wire seg_10_19_sp4_h_r_22_39808;
  wire seg_10_19_sp4_r_v_b_15_43405;
  wire seg_10_19_sp4_r_v_b_3_43281;
  wire seg_10_19_sp4_r_v_b_7_43285;
  wire seg_10_19_sp4_v_b_15_39574;
  wire seg_10_19_sp4_v_b_17_39576;
  wire seg_10_1_glb_netwk_0_5;
  wire seg_10_1_glb_netwk_4_9;
  wire seg_10_1_local_g0_1_41289;
  wire seg_10_1_local_g0_4_41292;
  wire seg_10_1_local_g0_5_41293;
  wire seg_10_1_local_g0_6_41294;
  wire seg_10_1_local_g1_3_41299;
  wire seg_10_1_local_g1_6_41302;
  wire seg_10_1_local_g1_7_41303;
  wire seg_10_1_local_g2_5_41309;
  wire seg_10_1_lutff_1_out_37416;
  wire seg_10_1_lutff_2_out_37417;
  wire seg_10_1_lutff_5_out_37420;
  wire seg_10_1_lutff_6_out_37421;
  wire seg_10_1_lutff_7_out_37422;
  wire seg_10_1_neigh_op_lft_1_33585;
  wire seg_10_1_neigh_op_lft_3_33587;
  wire seg_10_1_neigh_op_lft_4_33588;
  wire seg_10_1_neigh_op_lft_6_33590;
  wire seg_10_1_neigh_op_top_5_37548;
  wire seg_10_1_neigh_op_top_7_37550;
  wire seg_10_1_sp4_h_r_1_41387;
  wire seg_10_1_sp4_h_r_9_41397;
  wire seg_10_1_sp4_r_v_b_47_41440;
  wire seg_10_21_sp4_v_b_0_39695;
  wire seg_10_21_sp4_v_b_7_39700;
  wire seg_10_25_sp4_v_b_7_40192;
  wire seg_10_25_sp4_v_b_8_40195;
  wire seg_10_29_sp4_v_b_3_40680;
  wire seg_10_2_glb_netwk_0_5;
  wire seg_10_2_glb_netwk_4_9;
  wire seg_10_2_local_g0_1_41452;
  wire seg_10_2_local_g0_6_41457;
  wire seg_10_2_local_g0_7_41458;
  wire seg_10_2_local_g2_3_41470;
  wire seg_10_2_local_g2_7_41474;
  wire seg_10_2_local_g3_0_41475;
  wire seg_10_2_local_g3_2_41477;
  wire seg_10_2_local_g3_4_41479;
  wire seg_10_2_lutff_0_out_37543;
  wire seg_10_2_lutff_1_out_37544;
  wire seg_10_2_lutff_2_out_37545;
  wire seg_10_2_lutff_3_out_37546;
  wire seg_10_2_lutff_4_out_37547;
  wire seg_10_2_lutff_5_out_37548;
  wire seg_10_2_lutff_6_out_37549;
  wire seg_10_2_lutff_7_out_37550;
  wire seg_10_2_sp4_h_r_28_33889;
  wire seg_10_2_sp4_h_r_9_41556;
  wire seg_10_2_sp4_v_b_23_37595;
  wire seg_10_2_sp4_v_b_39_37729;
  wire seg_10_2_sp4_v_t_44_37857;
  wire seg_10_3_glb_netwk_0_5;
  wire seg_10_3_glb_netwk_4_9;
  wire seg_10_3_local_g1_2_41584;
  wire seg_10_3_local_g1_7_41589;
  wire seg_10_3_local_g2_3_41593;
  wire seg_10_3_local_g2_4_41594;
  wire seg_10_3_local_g2_5_41595;
  wire seg_10_3_local_g3_0_41598;
  wire seg_10_3_local_g3_5_41603;
  wire seg_10_3_local_g3_6_41604;
  wire seg_10_3_lutff_0_out_37702;
  wire seg_10_3_lutff_1_out_37703;
  wire seg_10_3_lutff_2_out_37704;
  wire seg_10_3_lutff_3_out_37705;
  wire seg_10_3_lutff_4_out_37706;
  wire seg_10_3_lutff_5_out_37707;
  wire seg_10_3_lutff_6_out_37708;
  wire seg_10_3_lutff_7_out_37709;
  wire seg_10_3_sp4_h_l_46_26914;
  wire seg_10_3_sp4_h_r_0_41668;
  wire seg_10_3_sp4_h_r_23_37839;
  wire seg_10_3_sp4_h_r_27_34011;
  wire seg_10_3_sp4_h_r_2_41672;
  wire seg_10_3_sp4_h_r_37_30175;
  wire seg_10_3_sp4_h_r_45_30185;
  wire seg_10_3_sp4_r_v_b_16_41433;
  wire seg_10_3_sp4_r_v_b_22_41439;
  wire seg_10_3_sp4_v_b_12_37597;
  wire seg_10_3_sp4_v_b_36_37849;
  wire seg_10_3_sp4_v_t_47_37983;
  wire seg_10_4_glb_netwk_0_5;
  wire seg_10_4_glb_netwk_3_8;
  wire seg_10_4_local_g0_6_41703;
  wire seg_10_4_local_g0_7_41704;
  wire seg_10_4_local_g1_1_41706;
  wire seg_10_4_local_g1_3_41708;
  wire seg_10_4_local_g1_5_41710;
  wire seg_10_4_local_g1_7_41712;
  wire seg_10_4_local_g2_1_41714;
  wire seg_10_4_local_g2_6_41719;
  wire seg_10_4_local_g3_3_41724;
  wire seg_10_4_local_g3_4_41725;
  wire seg_10_4_local_g3_6_41727;
  wire seg_10_4_lutff_1_out_37826;
  wire seg_10_4_lutff_3_out_37828;
  wire seg_10_4_lutff_6_out_37831;
  wire seg_10_4_neigh_op_lft_6_34000;
  wire seg_10_4_neigh_op_lft_7_34001;
  wire seg_10_4_sp12_v_b_16_41270;
  wire seg_10_4_sp4_h_r_10_41793;
  wire seg_10_4_sp4_h_r_19_37968;
  wire seg_10_4_sp4_h_r_1_41792;
  wire seg_10_4_sp4_h_r_23_37962;
  wire seg_10_4_sp4_h_r_27_34134;
  wire seg_10_4_sp4_h_r_30_34137;
  wire seg_10_4_sp4_h_r_3_41796;
  wire seg_10_4_sp4_h_r_5_41798;
  wire seg_10_4_sp4_r_v_b_31_41686;
  wire seg_10_4_sp4_v_b_1_37597;
  wire seg_10_4_sp4_v_b_36_37972;
  wire seg_10_4_sp4_v_t_37_38096;
  wire seg_10_4_sp4_v_t_41_38100;
  wire seg_10_5_glb_netwk_0_5;
  wire seg_10_5_glb_netwk_4_9;
  wire seg_10_5_local_g1_0_41828;
  wire seg_10_5_local_g1_4_41832;
  wire seg_10_5_local_g2_6_41842;
  wire seg_10_5_local_g3_2_41846;
  wire seg_10_5_local_g3_5_41849;
  wire seg_10_5_lutff_4_out_37952;
  wire seg_10_5_lutff_5_out_37953;
  wire seg_10_5_lutff_7_out_37955;
  wire seg_10_5_neigh_op_lft_0_34117;
  wire seg_10_5_neigh_op_tnl_2_34242;
  wire seg_10_5_sp4_r_v_b_38_41928;
  wire seg_10_5_sp4_v_b_12_37849;
  wire seg_10_5_sp4_v_b_2_37729;
  wire seg_10_5_sp4_v_b_9_37734;
  wire seg_10_6_glb_netwk_0_5;
  wire seg_10_6_glb_netwk_5_10;
  wire seg_10_6_local_g1_2_41953;
  wire seg_10_6_local_g2_1_41960;
  wire seg_10_6_local_g3_1_41968;
  wire seg_10_6_neigh_op_bnr_2_41781;
  wire seg_10_6_neigh_op_rgt_1_41903;
  wire seg_10_6_sp4_h_r_24_34375;
  wire seg_10_6_sp4_h_r_2_42041;
  wire seg_10_6_sp4_h_r_8_42047;
  wire seg_10_6_sp4_v_b_25_38095;
  wire seg_10_6_sp4_v_b_30_38102;
  wire seg_10_6_sp4_v_t_42_38347;
  wire seg_10_7_glb_netwk_0_5;
  wire seg_10_7_glb_netwk_4_9;
  wire seg_10_7_local_g0_4_42070;
  wire seg_10_7_local_g0_6_42072;
  wire seg_10_7_local_g0_7_42073;
  wire seg_10_7_local_g1_0_42074;
  wire seg_10_7_local_g2_0_42082;
  wire seg_10_7_local_g3_1_42091;
  wire seg_10_7_local_g3_3_42093;
  wire seg_10_7_lutff_0_out_38194;
  wire seg_10_7_lutff_1_out_38195;
  wire seg_10_7_lutff_3_out_38197;
  wire seg_10_7_lutff_7_out_38201;
  wire seg_10_7_neigh_op_lft_0_34363;
  wire seg_10_7_neigh_op_tnl_3_34489;
  wire seg_10_7_neigh_op_top_4_38321;
  wire seg_10_7_sp12_h_r_0_42156;
  wire seg_10_7_sp4_h_r_16_38336;
  wire seg_10_7_sp4_h_r_24_34498;
  wire seg_10_7_sp4_h_r_5_42167;
  wire seg_10_7_sp4_r_v_b_33_42057;
  wire seg_10_7_sp4_r_v_b_8_41812;
  wire seg_10_7_sp4_v_b_10_37983;
  wire seg_10_7_sp4_v_b_24_38219;
  wire seg_10_7_sp4_v_b_3_37974;
  wire seg_10_7_sp4_v_b_41_38346;
  wire seg_10_7_sp4_v_b_6_37979;
  wire seg_10_7_sp4_v_t_36_38464;
  wire seg_10_8_glb_netwk_0_5;
  wire seg_10_8_glb_netwk_4_9;
  wire seg_10_8_local_g0_4_42193;
  wire seg_10_8_local_g1_1_42198;
  wire seg_10_8_local_g1_2_42199;
  wire seg_10_8_local_g1_5_42202;
  wire seg_10_8_local_g1_6_42203;
  wire seg_10_8_local_g3_0_42213;
  wire seg_10_8_local_g3_5_42218;
  wire seg_10_8_lutff_1_out_38318;
  wire seg_10_8_lutff_3_out_38320;
  wire seg_10_8_lutff_4_out_38321;
  wire seg_10_8_lutff_5_out_38322;
  wire seg_10_8_lutff_6_out_38323;
  wire seg_10_8_lutff_7_out_38324;
  wire seg_10_8_neigh_op_lft_2_34488;
  wire seg_10_8_neigh_op_lft_4_34490;
  wire seg_10_8_neigh_op_lft_5_34491;
  wire seg_10_8_neigh_op_lft_6_34492;
  wire seg_10_8_neigh_op_tnl_0_34609;
  wire seg_10_8_sp4_h_r_14_38457;
  wire seg_10_8_sp4_h_r_1_42284;
  wire seg_10_8_sp4_h_r_46_30793;
  wire seg_10_8_sp4_r_v_b_1_41926;
  wire seg_10_8_sp4_r_v_b_47_42306;
  wire seg_10_8_sp4_v_b_3_38097;
  wire seg_10_8_sp4_v_b_6_38102;
  wire seg_10_8_sp4_v_t_37_38588;
  wire seg_10_8_sp4_v_t_41_38592;
  wire seg_10_9_glb_netwk_0_5;
  wire seg_10_9_glb_netwk_5_10;
  wire seg_10_9_local_g0_7_42319;
  wire seg_10_9_neigh_op_bot_7_38324;
  wire seg_10_9_sp12_v_b_22_42281;
  wire seg_10_9_sp4_h_r_2_42410;
  wire seg_10_9_sp4_h_r_3_42411;
  wire seg_10_9_sp4_v_b_0_38219;
  wire seg_10_9_sp4_v_b_11_38228;
  wire seg_10_9_sp4_v_b_5_38222;
  wire seg_11_10_glb_netwk_0_5;
  wire seg_11_10_local_g0_2_46268;
  wire seg_11_10_local_g0_7_46273;
  wire seg_11_10_local_g2_1_46283;
  wire seg_11_10_local_g2_3_46285;
  wire seg_11_10_lutff_1_out_42395;
  wire seg_11_10_lutff_4_out_42398;
  wire seg_11_10_lutff_7_out_42401;
  wire seg_11_10_neigh_op_bot_7_42278;
  wire seg_11_10_neigh_op_rgt_1_46226;
  wire seg_11_10_sp4_h_l_36_31037;
  wire seg_11_10_sp4_h_l_42_31045;
  wire seg_11_10_sp4_h_l_44_31047;
  wire seg_11_10_sp4_h_r_3_46365;
  wire seg_11_10_sp4_h_r_7_46369;
  wire seg_11_10_sp4_h_r_8_46370;
  wire seg_11_10_sp4_r_v_b_33_46257;
  wire seg_11_10_sp4_v_b_35_42428;
  wire seg_11_11_glb_netwk_0_5;
  wire seg_11_11_glb_netwk_4_9;
  wire seg_11_11_local_g0_0_46389;
  wire seg_11_11_local_g0_3_46392;
  wire seg_11_11_local_g0_6_46395;
  wire seg_11_11_local_g1_0_46397;
  wire seg_11_11_local_g1_4_46401;
  wire seg_11_11_local_g1_5_46402;
  wire seg_11_11_local_g1_6_46403;
  wire seg_11_11_local_g2_0_46405;
  wire seg_11_11_local_g2_4_46409;
  wire seg_11_11_local_g2_5_46410;
  wire seg_11_11_local_g3_1_46414;
  wire seg_11_11_local_g3_4_46417;
  wire seg_11_11_lutff_1_out_42518;
  wire seg_11_11_lutff_4_out_42521;
  wire seg_11_11_lutff_5_out_42522;
  wire seg_11_11_lutff_6_out_42523;
  wire seg_11_11_neigh_op_bot_4_42398;
  wire seg_11_11_neigh_op_lft_6_38692;
  wire seg_11_11_sp12_h_r_22_2407;
  wire seg_11_11_sp12_v_b_22_46358;
  wire seg_11_11_sp12_v_b_4_45216;
  wire seg_11_11_sp4_h_l_38_31164;
  wire seg_11_11_sp4_h_l_41_31165;
  wire seg_11_11_sp4_h_r_16_42659;
  wire seg_11_11_sp4_h_r_24_38821;
  wire seg_11_11_sp4_h_r_2_46487;
  wire seg_11_11_sp4_h_r_3_46488;
  wire seg_11_11_sp4_h_r_7_46492;
  wire seg_11_11_sp4_r_v_b_0_46127;
  wire seg_11_11_sp4_r_v_b_15_46252;
  wire seg_11_11_sp4_r_v_b_21_46258;
  wire seg_11_11_sp4_r_v_b_23_46260;
  wire seg_11_11_sp4_r_v_b_44_46503;
  wire seg_11_11_sp4_r_v_b_5_46130;
  wire seg_11_11_sp4_v_b_0_42296;
  wire seg_11_11_sp4_v_b_10_42306;
  wire seg_11_11_sp4_v_b_11_42305;
  wire seg_11_11_sp4_v_b_1_42295;
  wire seg_11_11_sp4_v_b_6_42302;
  wire seg_11_11_sp4_v_t_38_42789;
  wire seg_11_12_glb_netwk_0_5;
  wire seg_11_12_glb_netwk_1_6;
  wire seg_11_12_glb_netwk_4_9;
  wire seg_11_12_local_g0_0_46512;
  wire seg_11_12_local_g0_6_46518;
  wire seg_11_12_local_g0_7_46519;
  wire seg_11_12_local_g1_2_46522;
  wire seg_11_12_local_g1_3_46523;
  wire seg_11_12_local_g1_7_46527;
  wire seg_11_12_local_g2_1_46529;
  wire seg_11_12_local_g2_2_46530;
  wire seg_11_12_local_g2_7_46535;
  wire seg_11_12_local_g3_0_46536;
  wire seg_11_12_local_g3_2_46538;
  wire seg_11_12_local_g3_4_46540;
  wire seg_11_12_local_g3_7_46543;
  wire seg_11_12_lutff_2_out_42642;
  wire seg_11_12_neigh_op_bnl_1_38687;
  wire seg_11_12_neigh_op_rgt_0_46471;
  wire seg_11_12_neigh_op_tnr_2_46596;
  wire seg_11_12_sp12_v_b_10_45743;
  wire seg_11_12_sp4_h_r_10_46608;
  wire seg_11_12_sp4_h_r_15_42779;
  wire seg_11_12_sp4_h_r_28_38950;
  wire seg_11_12_sp4_h_r_2_46610;
  wire seg_11_12_sp4_h_r_31_38953;
  wire seg_11_12_sp4_r_v_b_1_46249;
  wire seg_11_12_sp4_r_v_b_24_46496;
  wire seg_11_12_sp4_r_v_b_3_46251;
  wire seg_11_12_sp4_r_v_b_47_46629;
  wire seg_11_12_sp4_v_b_15_42544;
  wire seg_11_12_sp4_v_b_34_42675;
  wire seg_11_12_sp4_v_b_3_42420;
  wire seg_11_12_sp4_v_b_40_42791;
  wire seg_11_12_sp4_v_b_6_42425;
  wire seg_11_12_sp4_v_b_9_42426;
  wire seg_11_12_sp4_v_t_39_42913;
  wire seg_11_13_glb_netwk_0_5;
  wire seg_11_13_local_g0_1_46636;
  wire seg_11_13_local_g1_1_46644;
  wire seg_11_13_local_g2_2_46653;
  wire seg_11_13_local_g2_4_46655;
  wire seg_11_13_local_g3_1_46660;
  wire seg_11_13_local_g3_2_46661;
  wire seg_11_13_lutff_4_out_42767;
  wire seg_11_13_sp12_v_b_0_45216;
  wire seg_11_13_sp12_v_b_1_45215;
  wire seg_11_13_sp4_h_r_11_46732;
  wire seg_11_13_sp4_h_r_17_42904;
  wire seg_11_13_sp4_h_r_1_46730;
  wire seg_11_13_sp4_h_r_25_39068;
  wire seg_11_13_sp4_h_r_34_39069;
  wire seg_11_13_sp4_h_r_9_46740;
  wire seg_11_13_sp4_v_b_20_42672;
  wire seg_11_13_sp4_v_b_26_42790;
  wire seg_11_13_sp4_v_t_43_43040;
  wire seg_11_14_glb_netwk_0_5;
  wire seg_11_14_local_g0_0_46758;
  wire seg_11_14_local_g0_3_46761;
  wire seg_11_14_local_g0_4_46762;
  wire seg_11_14_local_g1_2_46768;
  wire seg_11_14_local_g1_5_46771;
  wire seg_11_14_local_g3_3_46785;
  wire seg_11_14_neigh_op_tnr_3_46843;
  wire seg_11_14_sp12_v_b_14_46235;
  wire seg_11_14_sp12_v_b_8_45867;
  wire seg_11_14_sp4_h_l_39_31532;
  wire seg_11_14_sp4_h_r_0_46852;
  wire seg_11_14_sp4_h_r_10_46854;
  wire seg_11_14_sp4_h_r_2_46856;
  wire seg_11_14_sp4_h_r_42_35368;
  wire seg_11_14_sp4_h_r_4_46858;
  wire seg_11_14_sp4_h_r_8_46862;
  wire seg_11_14_sp4_r_v_b_21_46627;
  wire seg_11_14_sp4_v_b_20_42795;
  wire seg_11_14_sp4_v_b_21_42796;
  wire seg_11_14_sp4_v_b_3_42666;
  wire seg_11_14_sp4_v_b_9_42672;
  wire seg_11_15_glb_netwk_0_5;
  wire seg_11_15_local_g0_1_46882;
  wire seg_11_15_local_g0_4_46885;
  wire seg_11_15_local_g0_6_46887;
  wire seg_11_15_local_g1_7_46896;
  wire seg_11_15_local_g2_0_46897;
  wire seg_11_15_local_g2_2_46899;
  wire seg_11_15_local_g2_4_46901;
  wire seg_11_15_local_g2_5_46902;
  wire seg_11_15_local_g2_7_46904;
  wire seg_11_15_local_g3_5_46910;
  wire seg_11_15_local_g3_6_46911;
  wire seg_11_15_lutff_0_out_43009;
  wire seg_11_15_lutff_6_out_43015;
  wire seg_11_15_neigh_op_rgt_2_46842;
  wire seg_11_15_sp4_h_l_36_31652;
  wire seg_11_15_sp4_h_r_0_46975;
  wire seg_11_15_sp4_h_r_30_39321;
  wire seg_11_15_sp4_h_r_46_35485;
  wire seg_11_15_sp4_h_r_9_46986;
  wire seg_11_15_sp4_r_v_b_12_46741;
  wire seg_11_15_sp4_r_v_b_13_46742;
  wire seg_11_15_sp4_r_v_b_21_46750;
  wire seg_11_15_sp4_v_b_10_42798;
  wire seg_11_15_sp4_v_b_11_42797;
  wire seg_11_15_sp4_v_b_17_42915;
  wire seg_11_15_sp4_v_b_1_42787;
  wire seg_11_15_sp4_v_b_20_42918;
  wire seg_11_15_sp4_v_b_24_43034;
  wire seg_11_15_sp4_v_b_34_43044;
  wire seg_11_15_sp4_v_b_36_43156;
  wire seg_11_15_sp4_v_b_39_43159;
  wire seg_11_15_sp4_v_b_5_42791;
  wire seg_11_15_sp4_v_b_6_42794;
  wire seg_11_15_sp4_v_b_7_42793;
  wire seg_11_15_sp4_v_t_38_43281;
  wire seg_11_16_glb_netwk_0_5;
  wire seg_11_16_glb_netwk_1_6;
  wire seg_11_16_glb_netwk_4_9;
  wire seg_11_16_local_g0_4_47008;
  wire seg_11_16_local_g1_0_47012;
  wire seg_11_16_local_g1_1_47013;
  wire seg_11_16_local_g1_6_47018;
  wire seg_11_16_local_g2_2_47022;
  wire seg_11_16_local_g2_3_47023;
  wire seg_11_16_local_g3_2_47030;
  wire seg_11_16_local_g3_3_47031;
  wire seg_11_16_local_g3_5_47033;
  wire seg_11_16_lutff_3_out_43135;
  wire seg_11_16_lutff_4_out_43136;
  wire seg_11_16_sp12_v_b_2_45743;
  wire seg_11_16_sp4_h_l_40_31781;
  wire seg_11_16_sp4_h_r_17_43273;
  wire seg_11_16_sp4_h_r_18_43276;
  wire seg_11_16_sp4_h_r_22_43270;
  wire seg_11_16_sp4_h_r_26_39440;
  wire seg_11_16_sp4_h_r_27_39441;
  wire seg_11_16_sp4_r_v_b_45_47119;
  wire seg_11_16_sp4_v_b_32_43165;
  wire seg_11_16_sp4_v_b_6_42917;
  wire seg_11_16_sp4_v_b_8_42919;
  wire seg_11_16_sp4_v_t_39_43405;
  wire seg_11_17_glb_netwk_0_5;
  wire seg_11_17_local_g0_1_47128;
  wire seg_11_17_local_g0_2_47129;
  wire seg_11_17_local_g0_4_47131;
  wire seg_11_17_local_g0_5_47132;
  wire seg_11_17_local_g1_0_47135;
  wire seg_11_17_local_g1_1_47136;
  wire seg_11_17_local_g1_2_47137;
  wire seg_11_17_local_g1_3_47138;
  wire seg_11_17_local_g1_6_47141;
  wire seg_11_17_local_g2_0_47143;
  wire seg_11_17_local_g2_2_47145;
  wire seg_11_17_local_g3_5_47156;
  wire seg_11_17_lutff_0_out_43255;
  wire seg_11_17_lutff_2_out_43257;
  wire seg_11_17_lutff_3_out_43258;
  wire seg_11_17_lutff_4_out_43259;
  wire seg_11_17_lutff_5_out_43260;
  wire seg_11_17_lutff_6_out_43261;
  wire seg_11_17_lutff_7_out_43262;
  wire seg_11_17_sp12_v_b_5_45989;
  wire seg_11_17_sp4_h_r_12_43391;
  wire seg_11_17_sp4_h_r_13_43390;
  wire seg_11_17_sp4_h_r_1_47222;
  wire seg_11_17_sp4_h_r_22_43393;
  wire seg_11_17_sp4_h_r_6_47229;
  wire seg_11_17_sp4_r_v_b_10_46875;
  wire seg_11_17_sp4_r_v_b_1_46864;
  wire seg_11_17_sp4_v_b_0_43034;
  wire seg_11_17_sp4_v_b_10_43044;
  wire seg_11_17_sp4_v_b_3_43035;
  wire seg_11_18_glb_netwk_0_5;
  wire seg_11_18_local_g0_0_47250;
  wire seg_11_18_local_g0_1_47251;
  wire seg_11_18_local_g0_2_47252;
  wire seg_11_18_local_g0_5_47255;
  wire seg_11_18_local_g0_6_47256;
  wire seg_11_18_local_g0_7_47257;
  wire seg_11_18_local_g1_2_47260;
  wire seg_11_18_local_g1_5_47263;
  wire seg_11_18_local_g1_6_47264;
  wire seg_11_18_local_g1_7_47265;
  wire seg_11_18_local_g2_0_47266;
  wire seg_11_18_local_g2_2_47268;
  wire seg_11_18_local_g3_3_47277;
  wire seg_11_18_local_g3_4_47278;
  wire seg_11_18_local_g3_6_47280;
  wire seg_11_18_lutff_1_out_43379;
  wire seg_11_18_neigh_op_bot_5_43260;
  wire seg_11_18_neigh_op_bot_6_43261;
  wire seg_11_18_neigh_op_rgt_2_47211;
  wire seg_11_18_neigh_op_rgt_4_47213;
  wire seg_11_18_neigh_op_tnr_3_47335;
  wire seg_11_18_sp12_v_b_0_45867;
  wire seg_11_18_sp12_v_b_6_46235;
  wire seg_11_18_sp4_h_r_15_43517;
  wire seg_11_18_sp4_r_v_b_15_47113;
  wire seg_11_18_sp4_r_v_b_21_47119;
  wire seg_11_18_sp4_r_v_b_26_47236;
  wire seg_11_18_sp4_r_v_b_27_47235;
  wire seg_11_18_sp4_r_v_b_5_46991;
  wire seg_11_18_sp4_v_b_10_43167;
  wire seg_11_18_sp4_v_b_16_43283;
  wire seg_11_18_sp4_v_b_1_43156;
  wire seg_11_18_sp4_v_b_6_43163;
  wire seg_11_18_sp4_v_b_9_43164;
  wire seg_11_19_glb_netwk_0_5;
  wire seg_11_19_glb_netwk_7_12;
  wire seg_11_19_local_g1_1_47382;
  wire seg_11_19_lutff_1_out_43502;
  wire seg_11_19_sp4_v_b_9_43287;
  wire seg_11_1_glb_netwk_0_5;
  wire seg_11_1_glb_netwk_4_9;
  wire seg_11_1_local_g2_0_45135;
  wire seg_11_1_sp4_h_r_24_37555;
  wire seg_11_1_sp4_h_r_8_45227;
  wire seg_11_1_sp4_r_v_b_9_45276;
  wire seg_11_22_sp12_v_b_1_46358;
  wire seg_11_25_sp12_v_b_0_46728;
  wire seg_11_25_sp12_v_b_1_46727;
  wire seg_11_2_glb_netwk_0_5;
  wire seg_11_2_glb_netwk_4_9;
  wire seg_11_2_local_g0_1_45283;
  wire seg_11_2_local_g1_6_45296;
  wire seg_11_2_local_g2_1_45299;
  wire seg_11_2_local_g2_2_45300;
  wire seg_11_2_local_g2_3_45301;
  wire seg_11_2_local_g2_6_45304;
  wire seg_11_2_local_g2_7_45305;
  wire seg_11_2_local_g3_2_45308;
  wire seg_11_2_local_g3_5_45311;
  wire seg_11_2_local_g3_6_45312;
  wire seg_11_2_local_g3_7_45313;
  wire seg_11_2_lutff_2_out_41376;
  wire seg_11_2_lutff_4_out_41378;
  wire seg_11_2_lutff_7_out_41381;
  wire seg_11_2_neigh_op_bnl_1_37416;
  wire seg_11_2_neigh_op_bnl_2_37417;
  wire seg_11_2_neigh_op_bnl_7_37422;
  wire seg_11_2_neigh_op_bnr_1_45078;
  wire seg_11_2_neigh_op_rgt_3_45208;
  wire seg_11_2_sp4_h_r_10_45378;
  wire seg_11_2_sp4_h_r_11_45379;
  wire seg_11_2_sp4_h_r_1_45377;
  wire seg_11_2_sp4_h_r_22_41548;
  wire seg_11_2_sp4_h_r_28_37720;
  wire seg_11_2_sp4_h_r_34_37716;
  wire seg_11_2_sp4_h_r_4_45382;
  wire seg_11_2_sp4_v_b_26_41431;
  wire seg_11_2_sp4_v_b_30_41436;
  wire seg_11_2_sp4_v_b_37_41558;
  wire seg_11_2_sp4_v_b_38_41559;
  wire seg_11_2_sp4_v_b_39_41560;
  wire seg_11_3_local_g0_3_45408;
  wire seg_11_3_local_g0_6_45411;
  wire seg_11_3_local_g0_7_45412;
  wire seg_11_3_local_g1_0_45413;
  wire seg_11_3_local_g1_1_45414;
  wire seg_11_3_local_g1_2_45415;
  wire seg_11_3_local_g1_4_45417;
  wire seg_11_3_local_g1_5_45418;
  wire seg_11_3_local_g1_7_45420;
  wire seg_11_3_local_g2_4_45425;
  wire seg_11_3_local_g2_6_45427;
  wire seg_11_3_local_g3_0_45429;
  wire seg_11_3_local_g3_1_45430;
  wire seg_11_3_local_g3_6_45435;
  wire seg_11_3_lutff_1_out_41534;
  wire seg_11_3_lutff_2_out_41535;
  wire seg_11_3_lutff_3_out_41536;
  wire seg_11_3_lutff_4_out_41537;
  wire seg_11_3_lutff_5_out_41538;
  wire seg_11_3_lutff_6_out_41539;
  wire seg_11_3_lutff_7_out_41540;
  wire seg_11_3_neigh_op_bnl_1_37544;
  wire seg_11_3_neigh_op_bnl_4_37547;
  wire seg_11_3_neigh_op_bot_7_41381;
  wire seg_11_3_neigh_op_lft_0_37702;
  wire seg_11_3_neigh_op_lft_1_37703;
  wire seg_11_3_neigh_op_lft_2_37704;
  wire seg_11_3_neigh_op_lft_3_37705;
  wire seg_11_3_neigh_op_lft_4_37706;
  wire seg_11_3_neigh_op_lft_5_37707;
  wire seg_11_3_neigh_op_lft_6_37708;
  wire seg_11_3_neigh_op_lft_7_37709;
  wire seg_11_3_sp4_h_r_0_45499;
  wire seg_11_3_sp4_h_r_6_45507;
  wire seg_11_3_sp4_v_b_30_41564;
  wire seg_11_3_sp4_v_b_32_41566;
  wire seg_11_3_sp4_v_b_38_41682;
  wire seg_11_4_glb_netwk_0_5;
  wire seg_11_4_glb_netwk_4_9;
  wire seg_11_4_local_g0_1_45529;
  wire seg_11_4_local_g0_4_45532;
  wire seg_11_4_local_g0_5_45533;
  wire seg_11_4_local_g0_6_45534;
  wire seg_11_4_local_g1_2_45538;
  wire seg_11_4_local_g1_3_45539;
  wire seg_11_4_local_g1_5_45541;
  wire seg_11_4_local_g1_6_45542;
  wire seg_11_4_local_g1_7_45543;
  wire seg_11_4_local_g2_2_45546;
  wire seg_11_4_local_g3_2_45554;
  wire seg_11_4_local_g3_5_45557;
  wire seg_11_4_lutff_3_out_41659;
  wire seg_11_4_lutff_5_out_41661;
  wire seg_11_4_neigh_op_bot_1_41534;
  wire seg_11_4_neigh_op_bot_2_41535;
  wire seg_11_4_neigh_op_bot_3_41536;
  wire seg_11_4_neigh_op_bot_4_41537;
  wire seg_11_4_neigh_op_bot_5_41538;
  wire seg_11_4_neigh_op_bot_6_41539;
  wire seg_11_4_neigh_op_bot_7_41540;
  wire seg_11_4_neigh_op_rgt_5_45492;
  wire seg_11_4_sp12_h_r_6_34126;
  wire seg_11_4_sp4_h_l_40_30305;
  wire seg_11_4_sp4_h_l_46_30301;
  wire seg_11_4_sp4_h_r_0_45622;
  wire seg_11_4_sp4_h_r_1_45623;
  wire seg_11_4_sp4_h_r_26_37964;
  wire seg_11_4_sp4_h_r_28_37966;
  wire seg_11_4_sp4_h_r_3_45627;
  wire seg_11_4_sp4_h_r_5_45629;
  wire seg_11_4_sp4_h_r_6_45630;
  wire seg_11_4_sp4_h_r_7_45631;
  wire seg_11_4_sp4_h_r_8_45632;
  wire seg_11_4_sp4_r_v_b_5_45264;
  wire seg_11_4_sp4_v_b_10_41440;
  wire seg_11_4_sp4_v_b_14_41559;
  wire seg_11_4_sp4_v_b_2_41431;
  wire seg_11_4_sp4_v_t_36_41926;
  wire seg_11_4_sp4_v_t_37_41927;
  wire seg_11_4_sp4_v_t_40_41930;
  wire seg_11_4_sp4_v_t_41_41931;
  wire seg_11_5_glb_netwk_0_5;
  wire seg_11_5_glb_netwk_4_9;
  wire seg_11_5_local_g0_2_45653;
  wire seg_11_5_local_g0_3_45654;
  wire seg_11_5_local_g0_7_45658;
  wire seg_11_5_local_g1_3_45662;
  wire seg_11_5_local_g1_4_45663;
  wire seg_11_5_local_g1_6_45665;
  wire seg_11_5_local_g1_7_45666;
  wire seg_11_5_lutff_2_out_41781;
  wire seg_11_5_lutff_3_out_41782;
  wire seg_11_5_lutff_6_out_41785;
  wire seg_11_5_neigh_op_bot_3_41659;
  wire seg_11_5_neigh_op_lft_7_37955;
  wire seg_11_5_neigh_op_top_4_41906;
  wire seg_11_5_neigh_op_top_7_41909;
  wire seg_11_5_sp4_h_r_10_45747;
  wire seg_11_5_sp4_h_r_18_41923;
  wire seg_11_5_sp4_h_r_26_38087;
  wire seg_11_5_sp4_h_r_4_45751;
  wire seg_11_5_sp4_r_v_b_43_45764;
  wire seg_11_5_sp4_v_b_0_41558;
  wire seg_11_5_sp4_v_b_14_41682;
  wire seg_11_5_sp4_v_b_19_41687;
  wire seg_11_5_sp4_v_b_20_41688;
  wire seg_11_5_sp4_v_b_2_41560;
  wire seg_11_5_sp4_v_b_6_41564;
  wire seg_11_5_sp4_v_b_8_41566;
  wire seg_11_5_sp4_v_t_44_42057;
  wire seg_11_6_glb_netwk_0_5;
  wire seg_11_6_glb_netwk_4_9;
  wire seg_11_6_local_g2_0_45790;
  wire seg_11_6_local_g2_1_45791;
  wire seg_11_6_local_g2_3_45793;
  wire seg_11_6_local_g2_6_45796;
  wire seg_11_6_lutff_0_out_41902;
  wire seg_11_6_lutff_1_out_41903;
  wire seg_11_6_lutff_4_out_41906;
  wire seg_11_6_lutff_7_out_41909;
  wire seg_11_6_neigh_op_tnl_1_38195;
  wire seg_11_6_neigh_op_tnl_3_38197;
  wire seg_11_6_sp4_h_l_39_30548;
  wire seg_11_6_sp4_h_l_45_30554;
  wire seg_11_6_sp4_h_r_10_45870;
  wire seg_11_6_sp4_h_r_18_42046;
  wire seg_11_6_sp4_h_r_1_45869;
  wire seg_11_6_sp4_h_r_2_45872;
  wire seg_11_6_sp4_h_r_46_34378;
  wire seg_11_6_sp4_r_v_b_35_45767;
  wire seg_11_6_sp4_v_b_7_41686;
  wire seg_11_6_sp4_v_b_9_41688;
  wire seg_11_7_glb_netwk_0_5;
  wire seg_11_7_glb_netwk_5_10;
  wire seg_11_7_local_g1_0_45905;
  wire seg_11_7_local_g1_4_45909;
  wire seg_11_7_local_g3_2_45923;
  wire seg_11_7_neigh_op_lft_0_38194;
  wire seg_11_7_sp12_h_r_1_45988;
  wire seg_11_7_sp4_h_r_0_45991;
  wire seg_11_7_sp4_h_r_10_45993;
  wire seg_11_7_sp4_h_r_11_45994;
  wire seg_11_7_sp4_h_r_1_45992;
  wire seg_11_7_sp4_h_r_20_42171;
  wire seg_11_7_sp4_h_r_3_45996;
  wire seg_11_7_sp4_r_v_b_41_46008;
  wire seg_11_7_sp4_v_b_42_42178;
  wire seg_11_7_sp4_v_t_41_42300;
  wire seg_11_8_glb_netwk_0_5;
  wire seg_11_8_glb_netwk_4_9;
  wire seg_11_8_local_g0_1_46021;
  wire seg_11_8_local_g0_5_46025;
  wire seg_11_8_local_g1_0_46028;
  wire seg_11_8_local_g1_3_46031;
  wire seg_11_8_local_g1_5_46033;
  wire seg_11_8_local_g1_6_46034;
  wire seg_11_8_local_g2_4_46040;
  wire seg_11_8_local_g2_6_46042;
  wire seg_11_8_local_g2_7_46043;
  wire seg_11_8_lutff_0_out_42148;
  wire seg_11_8_lutff_1_out_42149;
  wire seg_11_8_lutff_2_out_42150;
  wire seg_11_8_lutff_4_out_42152;
  wire seg_11_8_neigh_op_lft_3_38320;
  wire seg_11_8_neigh_op_lft_6_38323;
  wire seg_11_8_sp12_h_r_14_19925;
  wire seg_11_8_sp12_h_r_20_7898;
  wire seg_11_8_sp12_h_r_22_1764;
  wire seg_11_8_sp12_v_b_10_45215;
  wire seg_11_8_sp4_h_l_38_30795;
  wire seg_11_8_sp4_h_l_43_30798;
  wire seg_11_8_sp4_h_l_46_30793;
  wire seg_11_8_sp4_h_r_0_46114;
  wire seg_11_8_sp4_h_r_11_46117;
  wire seg_11_8_sp4_h_r_16_42290;
  wire seg_11_8_sp4_h_r_20_42294;
  wire seg_11_8_sp4_h_r_21_42293;
  wire seg_11_8_sp4_h_r_38_34626;
  wire seg_11_8_sp4_h_r_3_46119;
  wire seg_11_8_sp4_h_r_42_34630;
  wire seg_11_8_sp4_h_r_44_34632;
  wire seg_11_8_sp4_h_r_46_34624;
  wire seg_11_8_sp4_h_r_5_46121;
  wire seg_11_8_sp4_r_v_b_14_45882;
  wire seg_11_8_sp4_r_v_b_15_45883;
  wire seg_11_8_sp4_r_v_b_17_45885;
  wire seg_11_8_sp4_r_v_b_21_45889;
  wire seg_11_8_sp4_r_v_b_33_46011;
  wire seg_11_8_sp4_v_b_4_41931;
  wire seg_11_8_sp4_v_b_7_41932;
  wire seg_11_9_glb_netwk_0_5;
  wire seg_11_9_glb_netwk_4_9;
  wire seg_11_9_local_g0_1_46144;
  wire seg_11_9_local_g1_3_46154;
  wire seg_11_9_local_g1_7_46158;
  wire seg_11_9_lutff_1_out_42272;
  wire seg_11_9_lutff_7_out_42278;
  wire seg_11_9_sp12_h_r_3_42402;
  wire seg_11_9_sp4_v_b_23_42183;
  wire seg_11_9_sp4_v_b_24_42296;
  wire seg_11_9_sp4_v_b_30_42302;
  wire seg_12_0_local_g0_5_48897;
  wire seg_12_0_local_g0_5_48897_i1;
  wire seg_12_0_local_g0_5_48897_i2;
  wire seg_12_0_local_g0_5_48897_i3;
  wire seg_12_0_logic_op_tnr_5_48913;
  wire seg_12_0_span4_vert_19_45240;
  wire seg_12_10_glb_netwk_0_5;
  wire seg_12_10_glb_netwk_4_9;
  wire seg_12_10_local_g0_0_50097;
  wire seg_12_10_local_g0_3_50100;
  wire seg_12_10_local_g0_4_50101;
  wire seg_12_10_local_g1_3_50108;
  wire seg_12_10_local_g1_5_50110;
  wire seg_12_10_local_g3_1_50122;
  wire seg_12_10_lutff_1_out_46226;
  wire seg_12_10_sp12_v_b_1_48926;
  wire seg_12_10_sp4_h_l_37_34867;
  wire seg_12_10_sp4_h_l_40_34874;
  wire seg_12_10_sp4_h_l_42_34876;
  wire seg_12_10_sp4_h_r_11_50194;
  wire seg_12_10_sp4_h_r_14_46365;
  wire seg_12_10_sp4_h_r_18_46369;
  wire seg_12_10_sp4_h_r_20_46371;
  wire seg_12_10_sp4_h_r_3_50196;
  wire seg_12_10_sp4_h_r_46_38701;
  wire seg_12_10_sp4_r_v_b_17_49962;
  wire seg_12_10_sp4_r_v_b_24_50081;
  wire seg_12_10_sp4_r_v_b_31_50086;
  wire seg_12_10_sp4_r_v_b_39_50206;
  wire seg_12_10_sp4_r_v_b_45_50212;
  wire seg_12_10_sp4_r_v_b_47_50214;
  wire seg_12_10_sp4_v_b_18_46132;
  wire seg_12_10_sp4_v_b_21_46135;
  wire seg_12_10_sp4_v_b_24_46250;
  wire seg_12_10_sp4_v_b_40_46376;
  wire seg_12_10_sp4_v_b_6_46010;
  wire seg_12_10_sp4_v_b_8_46012;
  wire seg_12_11_glb_netwk_0_5;
  wire seg_12_11_local_g0_2_50222;
  wire seg_12_11_local_g0_4_50224;
  wire seg_12_11_local_g0_7_50227;
  wire seg_12_11_local_g1_3_50231;
  wire seg_12_11_local_g1_5_50233;
  wire seg_12_11_local_g1_7_50235;
  wire seg_12_11_sp4_h_l_36_34991;
  wire seg_12_11_sp4_h_r_10_50316;
  wire seg_12_11_sp4_h_r_21_46493;
  wire seg_12_11_sp4_h_r_23_46485;
  wire seg_12_11_sp4_h_r_3_50319;
  wire seg_12_11_sp4_h_r_4_50320;
  wire seg_12_11_sp4_h_r_7_50323;
  wire seg_12_11_sp4_r_v_b_23_50091;
  wire seg_12_11_sp4_r_v_b_31_50209;
  wire seg_12_11_sp4_r_v_b_3_49959;
  wire seg_12_11_sp4_r_v_b_41_50331;
  wire seg_12_11_sp4_r_v_b_43_50333;
  wire seg_12_11_sp4_r_v_b_45_50335;
  wire seg_12_11_sp4_v_b_11_46136;
  wire seg_12_11_sp4_v_b_4_46131;
  wire seg_12_11_sp4_v_b_7_46132;
  wire seg_12_11_sp4_v_t_39_46621;
  wire seg_12_12_glb_netwk_0_5;
  wire seg_12_12_local_g0_2_50345;
  wire seg_12_12_local_g1_2_50353;
  wire seg_12_12_local_g1_4_50355;
  wire seg_12_12_local_g2_3_50362;
  wire seg_12_12_local_g2_4_50363;
  wire seg_12_12_local_g3_1_50368;
  wire seg_12_12_local_g3_5_50372;
  wire seg_12_12_lutff_0_out_46471;
  wire seg_12_12_lutff_1_out_46472;
  wire seg_12_12_neigh_op_rgt_5_50307;
  wire seg_12_12_neigh_op_top_2_46596;
  wire seg_12_12_sp12_v_b_0_48932;
  wire seg_12_12_sp4_h_l_38_35118;
  wire seg_12_12_sp4_h_l_46_35116;
  wire seg_12_12_sp4_h_r_10_50439;
  wire seg_12_12_sp4_h_r_12_46607;
  wire seg_12_12_sp4_h_r_2_50441;
  wire seg_12_12_sp4_h_r_6_50445;
  wire seg_12_12_sp4_r_v_b_35_50336;
  wire seg_12_12_sp4_v_b_0_46250;
  wire seg_12_12_sp4_v_b_10_46260;
  wire seg_12_12_sp4_v_b_2_46252;
  wire seg_12_12_sp4_v_b_44_46626;
  wire seg_12_12_sp4_v_b_4_46254;
  wire seg_12_12_sp4_v_b_8_46258;
  wire seg_12_12_sp4_v_t_38_46743;
  wire seg_12_12_sp4_v_t_42_46747;
  wire seg_12_12_sp4_v_t_44_46749;
  wire seg_12_13_glb_netwk_0_5;
  wire seg_12_13_glb_netwk_4_9;
  wire seg_12_13_local_g0_0_50466;
  wire seg_12_13_local_g0_6_50472;
  wire seg_12_13_local_g1_1_50475;
  wire seg_12_13_local_g1_2_50476;
  wire seg_12_13_local_g1_3_50477;
  wire seg_12_13_local_g3_2_50492;
  wire seg_12_13_local_g3_4_50494;
  wire seg_12_13_lutff_0_out_46594;
  wire seg_12_13_lutff_2_out_46596;
  wire seg_12_13_lutff_3_out_46597;
  wire seg_12_13_lutff_4_out_46598;
  wire seg_12_13_lutff_6_out_46600;
  wire seg_12_13_sp4_h_r_18_46738;
  wire seg_12_13_sp4_h_r_20_46740;
  wire seg_12_13_sp4_h_r_36_39068;
  wire seg_12_13_sp4_r_v_b_1_50203;
  wire seg_12_13_sp4_r_v_b_37_50573;
  wire seg_12_13_sp4_r_v_b_42_50578;
  wire seg_12_13_sp4_r_v_b_43_50579;
  wire seg_12_13_sp4_r_v_b_5_50207;
  wire seg_12_13_sp4_v_b_10_46383;
  wire seg_12_13_sp4_v_b_20_46503;
  wire seg_12_13_sp4_v_b_36_46741;
  wire seg_12_13_sp4_v_b_5_46376;
  wire seg_12_13_sp4_v_b_6_46379;
  wire seg_12_13_sp4_v_b_9_46380;
  wire seg_12_14_glb_netwk_0_5;
  wire seg_12_14_glb_netwk_1_6;
  wire seg_12_14_glb_netwk_4_9;
  wire seg_12_14_local_g0_1_50590;
  wire seg_12_14_local_g1_1_50598;
  wire seg_12_14_local_g1_2_50599;
  wire seg_12_14_local_g1_3_50600;
  wire seg_12_14_local_g1_5_50602;
  wire seg_12_14_local_g2_1_50606;
  wire seg_12_14_local_g2_4_50609;
  wire seg_12_14_local_g2_7_50612;
  wire seg_12_14_local_g3_1_50614;
  wire seg_12_14_local_g3_3_50616;
  wire seg_12_14_local_g3_4_50617;
  wire seg_12_14_local_g3_6_50619;
  wire seg_12_14_lutff_1_out_46718;
  wire seg_12_14_lutff_3_out_46720;
  wire seg_12_14_lutff_4_out_46721;
  wire seg_12_14_lutff_5_out_46722;
  wire seg_12_14_neigh_op_rgt_1_50549;
  wire seg_12_14_sp4_h_l_37_35359;
  wire seg_12_14_sp4_h_r_1_50684;
  wire seg_12_14_sp4_h_r_39_39194;
  wire seg_12_14_sp4_h_r_44_39201;
  wire seg_12_14_sp4_r_v_b_13_50450;
  wire seg_12_14_sp4_r_v_b_2_50329;
  wire seg_12_14_sp4_v_b_0_46496;
  wire seg_12_14_sp4_v_b_17_46623;
  wire seg_12_14_sp4_v_b_19_46625;
  wire seg_12_14_sp4_v_b_30_46748;
  wire seg_12_14_sp4_v_b_4_46500;
  wire seg_12_14_sp4_v_b_6_46502;
  wire seg_12_14_sp4_v_b_9_46503;
  wire seg_12_14_sp4_v_t_45_46996;
  wire seg_12_14_sp4_v_t_46_46997;
  wire seg_12_15_glb_netwk_0_5;
  wire seg_12_15_glb_netwk_4_9;
  wire seg_12_15_local_g0_2_50714;
  wire seg_12_15_local_g0_3_50715;
  wire seg_12_15_local_g1_3_50723;
  wire seg_12_15_local_g1_4_50724;
  wire seg_12_15_local_g2_3_50731;
  wire seg_12_15_local_g2_6_50734;
  wire seg_12_15_local_g3_3_50739;
  wire seg_12_15_local_g3_4_50740;
  wire seg_12_15_local_g3_6_50742;
  wire seg_12_15_lutff_0_out_46840;
  wire seg_12_15_lutff_2_out_46842;
  wire seg_12_15_lutff_3_out_46843;
  wire seg_12_15_lutff_4_out_46844;
  wire seg_12_15_lutff_5_out_46845;
  wire seg_12_15_neigh_op_bnr_2_50550;
  wire seg_12_15_neigh_op_tnr_3_50797;
  wire seg_12_15_neigh_op_top_3_46966;
  wire seg_12_15_sp4_h_l_37_35482;
  wire seg_12_15_sp4_h_l_41_35488;
  wire seg_12_15_sp4_h_r_0_50806;
  wire seg_12_15_sp4_h_r_12_46976;
  wire seg_12_15_sp4_h_r_20_46986;
  wire seg_12_15_sp4_h_r_22_46978;
  wire seg_12_15_sp4_h_r_30_43152;
  wire seg_12_15_sp4_h_r_34_43146;
  wire seg_12_15_sp4_h_r_36_39314;
  wire seg_12_15_sp4_h_r_38_39318;
  wire seg_12_15_sp4_h_r_4_50812;
  wire seg_12_15_sp4_r_v_b_15_50575;
  wire seg_12_15_sp4_r_v_b_19_50579;
  wire seg_12_15_sp4_r_v_b_21_50581;
  wire seg_12_15_sp4_r_v_b_23_50583;
  wire seg_12_15_sp4_r_v_b_31_50701;
  wire seg_12_15_sp4_r_v_b_3_50451;
  wire seg_12_15_sp4_r_v_b_5_50453;
  wire seg_12_15_sp4_r_v_b_7_50455;
  wire seg_12_15_sp4_v_b_14_46743;
  wire seg_12_15_sp4_v_b_18_46747;
  wire seg_12_15_sp4_v_b_20_46749;
  wire seg_12_15_sp4_v_b_2_46621;
  wire seg_12_15_sp4_v_b_34_46875;
  wire seg_12_15_sp4_v_b_36_46987;
  wire seg_12_15_sp4_v_b_38_46989;
  wire seg_12_15_sp4_v_b_3_46620;
  wire seg_12_15_sp4_v_b_46_46997;
  wire seg_12_15_sp4_v_b_8_46627;
  wire seg_12_15_sp4_v_t_39_47113;
  wire seg_12_16_glb_netwk_0_5;
  wire seg_12_16_glb_netwk_4_9;
  wire seg_12_16_local_g0_0_50835;
  wire seg_12_16_local_g0_1_50836;
  wire seg_12_16_local_g0_2_50837;
  wire seg_12_16_local_g0_3_50838;
  wire seg_12_16_local_g0_4_50839;
  wire seg_12_16_local_g0_5_50840;
  wire seg_12_16_local_g0_6_50841;
  wire seg_12_16_local_g0_7_50842;
  wire seg_12_16_local_g1_1_50844;
  wire seg_12_16_local_g1_3_50846;
  wire seg_12_16_local_g1_4_50847;
  wire seg_12_16_local_g1_5_50848;
  wire seg_12_16_local_g1_6_50849;
  wire seg_12_16_local_g1_7_50850;
  wire seg_12_16_local_g2_5_50856;
  wire seg_12_16_local_g2_6_50857;
  wire seg_12_16_local_g2_7_50858;
  wire seg_12_16_local_g3_5_50864;
  wire seg_12_16_local_g3_7_50866;
  wire seg_12_16_lutff_0_out_46963;
  wire seg_12_16_lutff_1_out_46964;
  wire seg_12_16_lutff_3_out_46966;
  wire seg_12_16_lutff_4_out_46967;
  wire seg_12_16_lutff_5_out_46968;
  wire seg_12_16_lutff_6_out_46969;
  wire seg_12_16_lutff_7_out_46970;
  wire seg_12_16_neigh_op_bot_5_46845;
  wire seg_12_16_neigh_op_rgt_7_50801;
  wire seg_12_16_neigh_op_tnr_5_50922;
  wire seg_12_16_neigh_op_tnr_7_50924;
  wire seg_12_16_neigh_op_top_1_47087;
  wire seg_12_16_neigh_op_top_2_47088;
  wire seg_12_16_neigh_op_top_3_47089;
  wire seg_12_16_neigh_op_top_6_47092;
  wire seg_12_16_neigh_op_top_7_47093;
  wire seg_12_16_sp12_v_b_4_49698;
  wire seg_12_16_sp4_h_r_11_50932;
  wire seg_12_16_sp4_h_r_16_47105;
  wire seg_12_16_sp4_h_r_29_43274;
  wire seg_12_16_sp4_h_r_4_50935;
  wire seg_12_16_sp4_r_v_b_6_50579;
  wire seg_12_16_sp4_v_b_10_46752;
  wire seg_12_16_sp4_v_b_11_46751;
  wire seg_12_16_sp4_v_b_1_46741;
  wire seg_12_16_sp4_v_b_20_46872;
  wire seg_12_16_sp4_v_b_4_46746;
  wire seg_12_16_sp4_v_b_8_46750;
  wire seg_12_16_sp4_v_b_9_46749;
  wire seg_12_16_sp4_v_t_38_47235;
  wire seg_12_17_glb_netwk_0_5;
  wire seg_12_17_glb_netwk_4_9;
  wire seg_12_17_local_g0_1_50959;
  wire seg_12_17_local_g1_0_50966;
  wire seg_12_17_local_g1_5_50971;
  wire seg_12_17_local_g2_4_50978;
  wire seg_12_17_lutff_1_out_47087;
  wire seg_12_17_lutff_2_out_47088;
  wire seg_12_17_lutff_3_out_47089;
  wire seg_12_17_lutff_4_out_47090;
  wire seg_12_17_lutff_6_out_47092;
  wire seg_12_17_lutff_7_out_47093;
  wire seg_12_17_neigh_op_bot_0_46963;
  wire seg_12_17_neigh_op_bot_1_46964;
  wire seg_12_17_neigh_op_bot_5_46968;
  wire seg_12_17_sp4_r_v_b_15_50821;
  wire seg_12_17_sp4_v_b_0_46865;
  wire seg_12_17_sp4_v_b_12_46987;
  wire seg_12_17_sp4_v_b_14_46989;
  wire seg_12_17_sp4_v_b_6_46871;
  wire seg_12_18_glb_netwk_0_5;
  wire seg_12_18_local_g0_1_51082;
  wire seg_12_18_local_g1_3_51092;
  wire seg_12_18_local_g1_4_51093;
  wire seg_12_18_lutff_2_out_47211;
  wire seg_12_18_lutff_4_out_47213;
  wire seg_12_18_sp4_h_r_3_51180;
  wire seg_12_18_sp4_r_v_b_25_51064;
  wire seg_12_18_sp4_v_b_11_46997;
  wire seg_12_18_sp4_v_b_4_46992;
  wire seg_12_19_glb_netwk_0_5;
  wire seg_12_19_local_g1_6_51218;
  wire seg_12_19_local_g3_3_51231;
  wire seg_12_19_lutff_3_out_47335;
  wire seg_12_19_sp4_r_v_b_19_51071;
  wire seg_12_19_sp4_v_b_22_47243;
  wire seg_12_1_glb_netwk_0_5;
  wire seg_12_1_glb_netwk_4_9;
  wire seg_12_1_local_g0_2_48952;
  wire seg_12_1_local_g0_4_48954;
  wire seg_12_1_local_g1_1_48959;
  wire seg_12_1_local_g2_1_48967;
  wire seg_12_1_local_g2_2_48968;
  wire seg_12_1_local_g3_1_48975;
  wire seg_12_1_local_g3_3_48977;
  wire seg_12_1_local_g3_5_48979;
  wire seg_12_1_lutff_1_out_45078;
  wire seg_12_1_lutff_2_out_45079;
  wire seg_12_1_lutff_3_out_45080;
  wire seg_12_1_lutff_4_out_45081;
  wire seg_12_1_neigh_op_tnr_1_49037;
  wire seg_12_1_sp4_h_r_11_49051;
  wire seg_12_1_sp4_h_r_42_37564;
  wire seg_12_1_sp4_r_v_b_19_49071;
  wire seg_12_1_sp4_r_v_b_21_49074;
  wire seg_12_1_sp4_r_v_b_23_49076;
  wire seg_12_1_sp4_r_v_b_25_49078;
  wire seg_12_1_sp4_r_v_b_35_49089;
  wire seg_12_1_sp4_r_v_b_37_49091;
  wire seg_12_1_sp4_r_v_b_39_49093;
  wire seg_12_1_sp4_r_v_b_41_49096;
  wire seg_12_1_sp4_r_v_b_45_49100;
  wire seg_12_1_sp4_v_b_34_45257;
  wire seg_12_1_sp4_v_b_9_45276;
  wire seg_12_22_sp12_v_b_1_50189;
  wire seg_12_2_glb_netwk_0_5;
  wire seg_12_2_glb_netwk_4_9;
  wire seg_12_2_local_g0_2_49115;
  wire seg_12_2_local_g0_6_49119;
  wire seg_12_2_local_g1_2_49123;
  wire seg_12_2_local_g1_3_49124;
  wire seg_12_2_local_g2_2_49131;
  wire seg_12_2_local_g2_5_49134;
  wire seg_12_2_lutff_0_out_45205;
  wire seg_12_2_lutff_2_out_45207;
  wire seg_12_2_lutff_3_out_45208;
  wire seg_12_2_lutff_6_out_45211;
  wire seg_12_2_neigh_op_bot_2_45079;
  wire seg_12_2_neigh_op_bot_3_45080;
  wire seg_12_2_neigh_op_lft_2_41376;
  wire seg_12_2_neigh_op_tnr_2_49197;
  wire seg_12_2_sp4_h_r_1_49208;
  wire seg_12_2_sp4_h_r_2_49211;
  wire seg_12_2_sp4_h_r_38_37719;
  wire seg_12_2_sp4_r_v_b_25_49090;
  wire seg_12_2_sp4_r_v_b_41_49224;
  wire seg_12_2_sp4_v_b_22_45258;
  wire seg_12_2_sp4_v_b_29_45264;
  wire seg_12_2_sp4_v_b_34_45271;
  wire seg_12_2_sp4_v_b_38_45390;
  wire seg_12_2_sp4_v_b_40_45392;
  wire seg_12_31_local_g1_6_52707;
  wire seg_12_31_local_g1_6_52707_i1;
  wire seg_12_31_local_g1_6_52707_i2;
  wire seg_12_31_local_g1_6_52707_i3;
  wire seg_12_31_span4_horz_r_6_48880;
  wire seg_12_3_glb_netwk_0_5;
  wire seg_12_3_glb_netwk_4_9;
  wire seg_12_3_local_g0_0_49236;
  wire seg_12_3_local_g0_2_49238;
  wire seg_12_3_local_g0_3_49239;
  wire seg_12_3_local_g0_4_49240;
  wire seg_12_3_local_g0_5_49241;
  wire seg_12_3_local_g1_2_49246;
  wire seg_12_3_local_g2_4_49256;
  wire seg_12_3_local_g2_5_49257;
  wire seg_12_3_local_g2_6_49258;
  wire seg_12_3_local_g3_6_49266;
  wire seg_12_3_lutff_4_out_45368;
  wire seg_12_3_lutff_5_out_45369;
  wire seg_12_3_lutff_6_out_45370;
  wire seg_12_3_neigh_op_bnl_4_41378;
  wire seg_12_3_neigh_op_bot_0_45205;
  wire seg_12_3_neigh_op_bot_2_45207;
  wire seg_12_3_neigh_op_rgt_6_49201;
  wire seg_12_3_neigh_op_tnl_5_41661;
  wire seg_12_3_neigh_op_tnr_6_49324;
  wire seg_12_3_neigh_op_top_3_45490;
  wire seg_12_3_sp12_v_b_14_48926;
  wire seg_12_3_sp4_h_l_42_34015;
  wire seg_12_3_sp4_h_l_43_34014;
  wire seg_12_3_sp4_h_r_24_41668;
  wire seg_12_3_sp4_h_r_28_41674;
  wire seg_12_3_sp4_h_r_40_37844;
  wire seg_12_3_sp4_h_r_8_49340;
  wire seg_12_3_sp4_r_v_b_25_49219;
  wire seg_12_3_sp4_r_v_b_45_49351;
  wire seg_12_3_sp4_v_b_10_45257;
  wire seg_12_3_sp4_v_b_11_45258;
  wire seg_12_3_sp4_v_b_12_45259;
  wire seg_12_3_sp4_v_b_24_45389;
  wire seg_12_3_sp4_v_b_30_45395;
  wire seg_12_3_sp4_v_b_40_45515;
  wire seg_12_4_glb_netwk_0_5;
  wire seg_12_4_local_g0_4_49363;
  wire seg_12_4_local_g0_6_49365;
  wire seg_12_4_local_g0_7_49366;
  wire seg_12_4_local_g1_0_49367;
  wire seg_12_4_local_g1_4_49371;
  wire seg_12_4_local_g1_6_49373;
  wire seg_12_4_local_g2_0_49375;
  wire seg_12_4_local_g2_3_49378;
  wire seg_12_4_local_g2_4_49379;
  wire seg_12_4_local_g2_5_49380;
  wire seg_12_4_local_g3_0_49383;
  wire seg_12_4_local_g3_1_49384;
  wire seg_12_4_local_g3_2_49385;
  wire seg_12_4_local_g3_3_49386;
  wire seg_12_4_local_g3_5_49388;
  wire seg_12_4_local_g3_7_49390;
  wire seg_12_4_lutff_0_out_45487;
  wire seg_12_4_lutff_3_out_45490;
  wire seg_12_4_lutff_4_out_45491;
  wire seg_12_4_lutff_5_out_45492;
  wire seg_12_4_neigh_op_bot_4_45368;
  wire seg_12_4_neigh_op_bot_6_45370;
  wire seg_12_4_neigh_op_rgt_0_49318;
  wire seg_12_4_neigh_op_rgt_3_49321;
  wire seg_12_4_neigh_op_tnl_3_41782;
  wire seg_12_4_sp4_h_r_10_49455;
  wire seg_12_4_sp4_h_r_11_49456;
  wire seg_12_4_sp4_h_r_14_45627;
  wire seg_12_4_sp4_h_r_18_45631;
  wire seg_12_4_sp4_h_r_23_45624;
  wire seg_12_4_sp4_h_r_29_41798;
  wire seg_12_4_sp4_h_r_31_41800;
  wire seg_12_4_sp4_h_r_33_41802;
  wire seg_12_4_sp4_h_r_34_41793;
  wire seg_12_4_sp4_h_r_5_49460;
  wire seg_12_4_sp4_h_r_6_49461;
  wire seg_12_4_sp4_h_r_9_49464;
  wire seg_12_4_sp4_r_v_b_29_49346;
  wire seg_12_4_sp4_r_v_b_4_49096;
  wire seg_12_4_sp4_v_b_10_45271;
  wire seg_12_4_sp4_v_b_1_45259;
  wire seg_12_4_sp4_v_b_32_45520;
  wire seg_12_4_sp4_v_b_36_45634;
  wire seg_12_4_sp4_v_t_46_45767;
  wire seg_12_5_glb_netwk_0_5;
  wire seg_12_5_glb_netwk_7_12;
  wire seg_12_5_local_g1_3_49493;
  wire seg_12_5_local_g1_4_49494;
  wire seg_12_5_local_g1_5_49495;
  wire seg_12_5_local_g3_5_49511;
  wire seg_12_5_neigh_op_bnr_4_49322;
  wire seg_12_5_sp4_h_r_0_49576;
  wire seg_12_5_sp4_h_r_10_49578;
  wire seg_12_5_sp4_r_v_b_13_49343;
  wire seg_12_5_sp4_r_v_b_21_49351;
  wire seg_12_5_sp4_v_b_0_45389;
  wire seg_12_5_sp4_v_b_36_45757;
  wire seg_12_5_sp4_v_b_3_45390;
  wire seg_12_5_sp4_v_b_5_45392;
  wire seg_12_5_sp4_v_b_6_45395;
  wire seg_12_5_sp4_v_t_41_45885;
  wire seg_12_5_sp4_v_t_45_45889;
  wire seg_12_6_glb_netwk_0_5;
  wire seg_12_6_glb_netwk_4_9;
  wire seg_12_6_local_g0_3_49608;
  wire seg_12_6_local_g0_5_49610;
  wire seg_12_6_local_g1_3_49616;
  wire seg_12_6_local_g1_4_49617;
  wire seg_12_6_local_g1_7_49620;
  wire seg_12_6_local_g2_2_49623;
  wire seg_12_6_local_g3_0_49629;
  wire seg_12_6_local_g3_1_49630;
  wire seg_12_6_local_g3_7_49636;
  wire seg_12_6_lutff_0_out_45733;
  wire seg_12_6_lutff_1_out_45734;
  wire seg_12_6_lutff_2_out_45735;
  wire seg_12_6_lutff_3_out_45736;
  wire seg_12_6_lutff_7_out_45740;
  wire seg_12_6_sp12_v_b_12_48932;
  wire seg_12_6_sp12_v_t_23_49698;
  wire seg_12_6_sp4_h_l_37_34375;
  wire seg_12_6_sp4_h_r_11_49702;
  wire seg_12_6_sp4_h_r_20_45879;
  wire seg_12_6_sp4_h_r_3_49704;
  wire seg_12_6_sp4_h_r_40_38213;
  wire seg_12_6_sp4_h_r_6_49707;
  wire seg_12_6_sp4_h_r_7_49708;
  wire seg_12_6_sp4_v_b_40_45884;
  wire seg_12_6_sp4_v_b_42_45886;
  wire seg_12_6_sp4_v_b_44_45888;
  wire seg_12_6_sp4_v_b_5_45515;
  wire seg_12_6_sp4_v_t_41_46008;
  wire seg_12_6_sp4_v_t_44_46011;
  wire seg_12_7_glb_netwk_0_5;
  wire seg_12_7_glb_netwk_3_8;
  wire seg_12_7_local_g1_1_49737;
  wire seg_12_7_local_g1_3_49739;
  wire seg_12_7_local_g1_5_49741;
  wire seg_12_7_local_g1_6_49742;
  wire seg_12_7_local_g2_0_49744;
  wire seg_12_7_local_g2_1_49745;
  wire seg_12_7_local_g2_6_49750;
  wire seg_12_7_local_g3_0_49752;
  wire seg_12_7_local_g3_3_49755;
  wire seg_12_7_lutff_0_out_45856;
  wire seg_12_7_lutff_1_out_45857;
  wire seg_12_7_lutff_6_out_45862;
  wire seg_12_7_lutff_7_out_45863;
  wire seg_12_7_neigh_op_tnl_0_42148;
  wire seg_12_7_sp4_h_r_22_45994;
  wire seg_12_7_sp4_h_r_24_42160;
  wire seg_12_7_sp4_h_r_25_42161;
  wire seg_12_7_sp4_h_r_2_49826;
  wire seg_12_7_sp4_h_r_40_38336;
  wire seg_12_7_sp4_h_r_4_49828;
  wire seg_12_7_sp4_r_v_b_14_49590;
  wire seg_12_7_sp4_r_v_b_19_49595;
  wire seg_12_7_sp4_r_v_b_5_49469;
  wire seg_12_7_sp4_v_b_19_45764;
  wire seg_12_7_sp4_v_b_1_45634;
  wire seg_12_7_sp4_v_b_2_45637;
  wire seg_12_7_sp4_v_t_36_46126;
  wire seg_12_8_glb_netwk_0_5;
  wire seg_12_8_glb_netwk_5_10;
  wire seg_12_8_local_g0_4_49855;
  wire seg_12_8_local_g0_6_49857;
  wire seg_12_8_local_g1_0_49859;
  wire seg_12_8_local_g1_2_49861;
  wire seg_12_8_neigh_op_lft_0_42148;
  wire seg_12_8_neigh_op_lft_2_42150;
  wire seg_12_8_sp4_h_r_0_49945;
  wire seg_12_8_sp4_h_r_4_49951;
  wire seg_12_8_sp4_h_r_5_49952;
  wire seg_12_8_sp4_h_r_8_49955;
  wire seg_12_8_sp4_h_r_9_49956;
  wire seg_12_8_sp4_r_v_b_27_49836;
  wire seg_12_8_sp4_v_b_12_45880;
  wire seg_12_8_sp4_v_b_1_45757;
  wire seg_12_8_sp4_v_b_46_46136;
  wire seg_12_8_sp4_v_b_6_45764;
  wire seg_12_8_sp4_v_t_36_46249;
  wire seg_12_9_glb_netwk_0_5;
  wire seg_12_9_local_g1_3_49985;
  wire seg_12_9_local_g2_3_49993;
  wire seg_12_9_local_g3_0_49998;
  wire seg_12_9_local_g3_3_50001;
  wire seg_12_9_sp4_h_r_28_42412;
  wire seg_12_9_sp4_h_r_2_50072;
  wire seg_12_9_sp4_h_r_32_42416;
  wire seg_12_9_sp4_h_r_3_50073;
  wire seg_12_9_sp4_r_v_b_11_49721;
  wire seg_12_9_sp4_r_v_b_43_50087;
  wire seg_12_9_sp4_v_b_3_45882;
  wire seg_12_9_sp4_v_b_40_46253;
  wire seg_12_9_sp4_v_b_43_46256;
  wire seg_12_9_sp4_v_b_5_45884;
  wire seg_12_9_sp4_v_b_6_45887;
  wire seg_12_9_sp4_v_b_7_45886;
  wire seg_12_9_sp4_v_b_9_45888;
  wire seg_13_0_local_g1_4_52735;
  wire seg_13_0_local_g1_4_52735_i1;
  wire seg_13_0_local_g1_4_52735_i2;
  wire seg_13_0_local_g1_4_52735_i3;
  wire seg_13_0_span4_horz_r_4_48940;
  wire seg_13_0_span4_vert_20_49073;
  wire seg_13_0_span4_vert_4_49094;
  wire seg_13_10_glb_netwk_0_5;
  wire seg_13_10_local_g0_1_53929;
  wire seg_13_10_local_g1_4_53940;
  wire seg_13_10_local_g1_5_53941;
  wire seg_13_10_local_g1_6_53942;
  wire seg_13_10_local_g2_0_53944;
  wire seg_13_10_local_g2_1_53945;
  wire seg_13_10_local_g2_2_53946;
  wire seg_13_10_local_g2_5_53949;
  wire seg_13_10_local_g3_0_53952;
  wire seg_13_10_local_g3_1_53953;
  wire seg_13_10_local_g3_3_53955;
  wire seg_13_10_lutff_1_out_50057;
  wire seg_13_10_lutff_2_out_50058;
  wire seg_13_10_lutff_5_out_50061;
  wire seg_13_10_sp12_v_b_16_53529;
  wire seg_13_10_sp4_h_l_44_38709;
  wire seg_13_10_sp4_h_l_47_38700;
  wire seg_13_10_sp4_h_r_4_54028;
  wire seg_13_10_sp4_h_r_8_54032;
  wire seg_13_10_sp4_r_v_b_25_53911;
  wire seg_13_10_sp4_r_v_b_34_53922;
  wire seg_13_10_sp4_r_v_b_37_54035;
  wire seg_13_10_sp4_r_v_b_6_53672;
  wire seg_13_10_sp4_r_v_b_9_53673;
  wire seg_13_10_sp4_v_b_21_49966;
  wire seg_13_10_sp4_v_b_35_50090;
  wire seg_13_10_sp4_v_b_40_50207;
  wire seg_13_10_sp4_v_b_6_49841;
  wire seg_13_10_sp4_v_t_46_50336;
  wire seg_13_11_glb_netwk_0_5;
  wire seg_13_11_local_g0_4_54055;
  wire seg_13_11_local_g0_5_54056;
  wire seg_13_11_local_g0_7_54058;
  wire seg_13_11_local_g1_7_54066;
  wire seg_13_11_local_g2_3_54070;
  wire seg_13_11_local_g2_5_54072;
  wire seg_13_11_local_g2_6_54073;
  wire seg_13_11_local_g3_3_54078;
  wire seg_13_11_local_g3_7_54082;
  wire seg_13_11_neigh_op_bot_5_50061;
  wire seg_13_11_neigh_op_top_4_50306;
  wire seg_13_11_sp12_v_b_18_53774;
  wire seg_13_11_sp12_v_b_20_53898;
  wire seg_13_11_sp4_h_l_38_38826;
  wire seg_13_11_sp4_h_l_40_38828;
  wire seg_13_11_sp4_h_l_47_38823;
  wire seg_13_11_sp4_h_r_23_50316;
  wire seg_13_11_sp4_h_r_2_54149;
  wire seg_13_11_sp4_h_r_4_54151;
  wire seg_13_11_sp4_h_r_5_54152;
  wire seg_13_11_sp4_h_r_8_54155;
  wire seg_13_11_sp4_r_v_b_11_53798;
  wire seg_13_11_sp4_v_b_10_49968;
  wire seg_13_11_sp4_v_b_1_49957;
  wire seg_13_11_sp4_v_b_27_50205;
  wire seg_13_11_sp4_v_b_29_50207;
  wire seg_13_11_sp4_v_b_31_50209;
  wire seg_13_11_sp4_v_b_44_50334;
  wire seg_13_11_sp4_v_b_46_50336;
  wire seg_13_11_sp4_v_b_7_49963;
  wire seg_13_11_sp4_v_t_37_50450;
  wire seg_13_11_sp4_v_t_38_50451;
  wire seg_13_11_sp4_v_t_40_50453;
  wire seg_13_11_sp4_v_t_42_50455;
  wire seg_13_11_sp4_v_t_43_50456;
  wire seg_13_12_glb_netwk_0_5;
  wire seg_13_12_local_g0_2_54176;
  wire seg_13_12_local_g0_5_54179;
  wire seg_13_12_local_g0_6_54180;
  wire seg_13_12_local_g1_1_54183;
  wire seg_13_12_local_g1_2_54184;
  wire seg_13_12_local_g2_5_54195;
  wire seg_13_12_local_g2_6_54196;
  wire seg_13_12_local_g3_1_54199;
  wire seg_13_12_local_g3_7_54205;
  wire seg_13_12_lutff_0_out_50302;
  wire seg_13_12_lutff_2_out_50304;
  wire seg_13_12_lutff_3_out_50305;
  wire seg_13_12_lutff_4_out_50306;
  wire seg_13_12_lutff_5_out_50307;
  wire seg_13_12_lutff_6_out_50308;
  wire seg_13_12_sp12_v_b_1_52762;
  wire seg_13_12_sp4_h_r_13_50437;
  wire seg_13_12_sp4_h_r_18_50446;
  wire seg_13_12_sp4_h_r_34_46608;
  wire seg_13_12_sp4_r_v_b_13_54035;
  wire seg_13_12_sp4_r_v_b_14_54036;
  wire seg_13_12_sp4_r_v_b_17_54039;
  wire seg_13_12_sp4_r_v_b_23_54045;
  wire seg_13_12_sp4_r_v_b_25_54157;
  wire seg_13_12_sp4_r_v_b_2_53914;
  wire seg_13_12_sp4_r_v_b_30_54164;
  wire seg_13_12_sp4_r_v_b_31_54163;
  wire seg_13_12_sp4_v_b_10_50091;
  wire seg_13_12_sp4_v_b_5_50084;
  wire seg_13_12_sp4_v_b_7_50086;
  wire seg_13_12_sp4_v_t_37_50573;
  wire seg_13_12_sp4_v_t_39_50575;
  wire seg_13_12_sp4_v_t_41_50577;
  wire seg_13_12_sp4_v_t_45_50581;
  wire seg_13_13_glb_netwk_0_5;
  wire seg_13_13_local_g0_2_54299;
  wire seg_13_13_local_g0_6_54303;
  wire seg_13_13_local_g0_7_54304;
  wire seg_13_13_local_g1_0_54305;
  wire seg_13_13_local_g1_2_54307;
  wire seg_13_13_local_g1_3_54308;
  wire seg_13_13_local_g1_4_54309;
  wire seg_13_13_local_g1_6_54311;
  wire seg_13_13_local_g2_0_54313;
  wire seg_13_13_local_g2_3_54316;
  wire seg_13_13_local_g2_4_54317;
  wire seg_13_13_local_g3_2_54323;
  wire seg_13_13_local_g3_3_54324;
  wire seg_13_13_local_g3_4_54325;
  wire seg_13_13_local_g3_5_54326;
  wire seg_13_13_lutff_0_out_50425;
  wire seg_13_13_lutff_2_out_50427;
  wire seg_13_13_lutff_3_out_50428;
  wire seg_13_13_lutff_5_out_50430;
  wire seg_13_13_neigh_op_bot_0_50302;
  wire seg_13_13_neigh_op_bot_2_50304;
  wire seg_13_13_neigh_op_bot_3_50305;
  wire seg_13_13_neigh_op_bot_6_50308;
  wire seg_13_13_neigh_op_lft_2_46596;
  wire seg_13_13_sp4_h_r_3_54396;
  wire seg_13_13_sp4_r_v_b_12_54157;
  wire seg_13_13_sp4_r_v_b_20_54165;
  wire seg_13_13_sp4_r_v_b_31_54286;
  wire seg_13_13_sp4_r_v_b_41_54408;
  wire seg_13_13_sp4_r_v_b_4_54039;
  wire seg_13_13_sp4_v_b_10_50214;
  wire seg_13_13_sp4_v_b_1_50203;
  wire seg_13_13_sp4_v_b_22_50336;
  wire seg_13_13_sp4_v_b_2_50206;
  wire seg_13_13_sp4_v_b_34_50460;
  wire seg_13_13_sp4_v_b_35_50459;
  wire seg_13_13_sp4_v_b_44_50580;
  wire seg_13_13_sp4_v_b_5_50207;
  wire seg_13_13_sp4_v_b_7_50209;
  wire seg_13_13_sp4_v_b_8_50212;
  wire seg_13_13_sp4_v_t_42_50701;
  wire seg_13_14_glb_netwk_0_5;
  wire seg_13_14_local_g0_5_54425;
  wire seg_13_14_local_g0_7_54427;
  wire seg_13_14_local_g1_0_54428;
  wire seg_13_14_local_g1_1_54429;
  wire seg_13_14_local_g1_3_54431;
  wire seg_13_14_local_g1_5_54433;
  wire seg_13_14_local_g1_7_54435;
  wire seg_13_14_local_g2_0_54436;
  wire seg_13_14_local_g2_1_54437;
  wire seg_13_14_local_g2_2_54438;
  wire seg_13_14_local_g3_0_54444;
  wire seg_13_14_local_g3_2_54446;
  wire seg_13_14_local_g3_3_54447;
  wire seg_13_14_local_g3_6_54450;
  wire seg_13_14_lutff_1_out_50549;
  wire seg_13_14_lutff_2_out_50550;
  wire seg_13_14_neigh_op_bnl_2_46596;
  wire seg_13_14_neigh_op_tnl_0_46840;
  wire seg_13_14_neigh_op_tnr_2_54504;
  wire seg_13_14_sp12_v_b_10_53651;
  wire seg_13_14_sp12_v_b_14_53897;
  wire seg_13_14_sp4_h_r_0_54514;
  wire seg_13_14_sp4_h_r_10_54516;
  wire seg_13_14_sp4_h_r_18_50692;
  wire seg_13_14_sp4_h_r_21_50693;
  wire seg_13_14_sp4_h_r_28_46858;
  wire seg_13_14_sp4_h_r_2_54518;
  wire seg_13_14_sp4_h_r_34_46854;
  wire seg_13_14_sp4_h_r_3_54519;
  wire seg_13_14_sp4_h_r_40_43028;
  wire seg_13_14_sp4_h_r_4_54520;
  wire seg_13_14_sp4_h_r_7_54523;
  wire seg_13_14_sp4_h_r_8_54524;
  wire seg_13_14_sp4_r_v_b_19_54287;
  wire seg_13_14_sp4_r_v_b_1_54157;
  wire seg_13_14_sp4_r_v_b_22_54290;
  wire seg_13_14_sp4_r_v_b_35_54413;
  wire seg_13_14_sp4_r_v_b_3_54159;
  wire seg_13_14_sp4_r_v_b_7_54163;
  wire seg_13_14_sp4_r_v_b_8_54166;
  wire seg_13_14_sp4_r_v_b_9_54165;
  wire seg_13_14_sp4_v_b_0_50327;
  wire seg_13_14_sp4_v_b_21_50458;
  wire seg_13_14_sp4_v_b_38_50697;
  wire seg_13_14_sp4_v_b_4_50331;
  wire seg_13_14_sp4_v_b_6_50333;
  wire seg_13_14_sp4_v_b_8_50335;
  wire seg_13_14_sp4_v_b_9_50334;
  wire seg_13_14_sp4_v_t_38_50820;
  wire seg_13_15_glb_netwk_0_5;
  wire seg_13_15_local_g0_0_54543;
  wire seg_13_15_local_g0_1_54544;
  wire seg_13_15_local_g0_3_54546;
  wire seg_13_15_local_g0_6_54549;
  wire seg_13_15_local_g1_0_54551;
  wire seg_13_15_local_g1_1_54552;
  wire seg_13_15_local_g1_2_54553;
  wire seg_13_15_local_g1_3_54554;
  wire seg_13_15_local_g1_4_54555;
  wire seg_13_15_local_g1_5_54556;
  wire seg_13_15_local_g2_2_54561;
  wire seg_13_15_local_g3_0_54567;
  wire seg_13_15_local_g3_7_54574;
  wire seg_13_15_lutff_1_out_50672;
  wire seg_13_15_lutff_2_out_50673;
  wire seg_13_15_neigh_op_bot_1_50549;
  wire seg_13_15_neigh_op_lft_3_46843;
  wire seg_13_15_neigh_op_lft_4_46844;
  wire seg_13_15_neigh_op_rgt_2_54504;
  wire seg_13_15_neigh_op_top_1_50795;
  wire seg_13_15_neigh_op_top_3_50797;
  wire seg_13_15_neigh_op_top_6_50800;
  wire seg_13_15_sp12_v_b_16_54144;
  wire seg_13_15_sp4_h_l_36_39314;
  wire seg_13_15_sp4_h_r_18_50815;
  wire seg_13_15_sp4_h_r_4_54643;
  wire seg_13_15_sp4_h_r_8_54647;
  wire seg_13_15_sp4_r_v_b_16_54407;
  wire seg_13_15_sp4_r_v_b_41_54654;
  wire seg_13_15_sp4_r_v_b_43_54656;
  wire seg_13_15_sp4_r_v_b_45_54658;
  wire seg_13_15_sp4_v_b_10_50460;
  wire seg_13_15_sp4_v_b_13_50573;
  wire seg_13_15_sp4_v_b_18_50578;
  wire seg_13_15_sp4_v_b_1_50449;
  wire seg_13_15_sp4_v_b_39_50821;
  wire seg_13_15_sp4_v_b_46_50828;
  wire seg_13_15_sp4_v_b_4_50454;
  wire seg_13_15_sp4_v_b_8_50458;
  wire seg_13_15_sp4_v_t_43_50948;
  wire seg_13_16_glb_netwk_0_5;
  wire seg_13_16_glb_netwk_4_9;
  wire seg_13_16_local_g0_1_54667;
  wire seg_13_16_local_g0_2_54668;
  wire seg_13_16_local_g0_3_54669;
  wire seg_13_16_local_g0_4_54670;
  wire seg_13_16_local_g0_6_54672;
  wire seg_13_16_local_g0_7_54673;
  wire seg_13_16_local_g1_2_54676;
  wire seg_13_16_local_g1_3_54677;
  wire seg_13_16_local_g1_4_54678;
  wire seg_13_16_local_g1_5_54679;
  wire seg_13_16_local_g2_0_54682;
  wire seg_13_16_local_g2_3_54685;
  wire seg_13_16_local_g3_4_54694;
  wire seg_13_16_local_g3_5_54695;
  wire seg_13_16_local_g3_6_54696;
  wire seg_13_16_lutff_1_out_50795;
  wire seg_13_16_lutff_2_out_50796;
  wire seg_13_16_lutff_3_out_50797;
  wire seg_13_16_lutff_4_out_50798;
  wire seg_13_16_lutff_5_out_50799;
  wire seg_13_16_lutff_6_out_50800;
  wire seg_13_16_lutff_7_out_50801;
  wire seg_13_16_neigh_op_bot_1_50672;
  wire seg_13_16_neigh_op_bot_2_50673;
  wire seg_13_16_neigh_op_lft_4_46967;
  wire seg_13_16_neigh_op_tnl_6_47092;
  wire seg_13_16_neigh_op_top_3_50920;
  wire seg_13_16_neigh_op_top_4_50921;
  wire seg_13_16_neigh_op_top_5_50922;
  wire seg_13_16_sp4_h_r_22_50932;
  wire seg_13_16_sp4_h_r_38_43272;
  wire seg_13_16_sp4_h_r_40_43274;
  wire seg_13_16_sp4_h_r_8_54770;
  wire seg_13_16_sp4_r_v_b_39_54775;
  wire seg_13_16_sp4_r_v_b_7_54409;
  wire seg_13_16_sp4_r_v_b_9_54411;
  wire seg_13_16_sp4_v_b_10_50583;
  wire seg_13_16_sp4_v_b_1_50572;
  wire seg_13_16_sp4_v_b_38_50943;
  wire seg_13_16_sp4_v_b_5_50576;
  wire seg_13_16_sp4_v_b_6_50579;
  wire seg_13_16_sp4_v_b_9_50580;
  wire seg_13_16_sp4_v_t_38_51066;
  wire seg_13_16_sp4_v_t_39_51067;
  wire seg_13_16_sp4_v_t_45_51073;
  wire seg_13_17_glb_netwk_0_5;
  wire seg_13_17_glb_netwk_4_9;
  wire seg_13_17_local_g0_0_54789;
  wire seg_13_17_local_g0_1_54790;
  wire seg_13_17_local_g0_4_54793;
  wire seg_13_17_local_g0_7_54796;
  wire seg_13_17_local_g1_3_54800;
  wire seg_13_17_local_g1_6_54803;
  wire seg_13_17_local_g1_7_54804;
  wire seg_13_17_local_g3_3_54816;
  wire seg_13_17_lutff_1_out_50918;
  wire seg_13_17_lutff_3_out_50920;
  wire seg_13_17_lutff_4_out_50921;
  wire seg_13_17_lutff_5_out_50922;
  wire seg_13_17_lutff_7_out_50924;
  wire seg_13_17_neigh_op_bot_3_50797;
  wire seg_13_17_neigh_op_lft_6_47092;
  wire seg_13_17_neigh_op_lft_7_47093;
  wire seg_13_17_sp4_h_r_11_54886;
  wire seg_13_17_sp4_h_r_14_51057;
  wire seg_13_17_sp4_h_r_30_47229;
  wire seg_13_17_sp4_h_r_46_43393;
  wire seg_13_17_sp4_r_v_b_15_54652;
  wire seg_13_17_sp4_v_b_14_50820;
  wire seg_13_17_sp4_v_b_30_50948;
  wire seg_13_17_sp4_v_b_3_50697;
  wire seg_13_17_sp4_v_b_7_50701;
  wire seg_13_17_sp4_v_b_8_50704;
  wire seg_13_18_glb_netwk_0_5;
  wire seg_13_18_local_g0_0_54912;
  wire seg_13_18_local_g0_1_54913;
  wire seg_13_18_local_g0_3_54915;
  wire seg_13_18_local_g0_4_54916;
  wire seg_13_18_local_g0_5_54917;
  wire seg_13_18_local_g0_7_54919;
  wire seg_13_18_local_g1_0_54920;
  wire seg_13_18_local_g1_3_54923;
  wire seg_13_18_local_g1_4_54924;
  wire seg_13_18_local_g1_5_54925;
  wire seg_13_18_local_g1_6_54926;
  wire seg_13_18_local_g1_7_54927;
  wire seg_13_18_local_g2_0_54928;
  wire seg_13_18_local_g2_1_54929;
  wire seg_13_18_local_g2_2_54930;
  wire seg_13_18_local_g2_3_54931;
  wire seg_13_18_local_g2_5_54933;
  wire seg_13_18_local_g2_7_54935;
  wire seg_13_18_local_g3_0_54936;
  wire seg_13_18_local_g3_2_54938;
  wire seg_13_18_local_g3_3_54939;
  wire seg_13_18_local_g3_5_54941;
  wire seg_13_18_local_g3_6_54942;
  wire seg_13_18_lutff_1_out_51041;
  wire seg_13_18_lutff_2_out_51042;
  wire seg_13_18_lutff_6_out_51046;
  wire seg_13_18_neigh_op_bot_7_50924;
  wire seg_13_18_sp12_v_b_0_53529;
  wire seg_13_18_sp12_v_b_2_53651;
  wire seg_13_18_sp12_v_b_5_53774;
  wire seg_13_18_sp12_v_b_6_53897;
  wire seg_13_18_sp12_v_b_7_53898;
  wire seg_13_18_sp4_h_r_14_51180;
  wire seg_13_18_sp4_h_r_25_47345;
  wire seg_13_18_sp4_h_r_38_43518;
  wire seg_13_18_sp4_r_v_b_18_54778;
  wire seg_13_18_sp4_r_v_b_19_54779;
  wire seg_13_18_sp4_r_v_b_24_54896;
  wire seg_13_18_sp4_r_v_b_27_54897;
  wire seg_13_18_sp4_r_v_b_4_54654;
  wire seg_13_18_sp4_r_v_b_5_54653;
  wire seg_13_18_sp4_r_v_b_6_54656;
  wire seg_13_18_sp4_r_v_b_8_54658;
  wire seg_13_18_sp4_v_b_10_50829;
  wire seg_13_18_sp4_v_b_11_50828;
  wire seg_13_18_sp4_v_b_26_51067;
  wire seg_13_18_sp4_v_b_29_51068;
  wire seg_13_18_sp4_v_b_32_51073;
  wire seg_13_18_sp4_v_b_3_50820;
  wire seg_13_18_sp4_v_b_43_51194;
  wire seg_13_18_sp4_v_b_4_50823;
  wire seg_13_18_sp4_v_b_5_50822;
  wire seg_13_18_sp4_v_b_6_50825;
  wire seg_13_18_sp4_v_b_7_50824;
  wire seg_13_18_sp4_v_b_8_50827;
  wire seg_13_18_sp4_v_b_9_50826;
  wire seg_13_19_glb_netwk_0_5;
  wire seg_13_19_local_g0_1_55036;
  wire seg_13_19_local_g0_4_55039;
  wire seg_13_19_local_g1_1_55044;
  wire seg_13_19_local_g1_3_55046;
  wire seg_13_19_local_g1_6_55049;
  wire seg_13_19_sp4_v_b_14_51066;
  wire seg_13_19_sp4_v_b_1_50941;
  wire seg_13_19_sp4_v_b_20_51072;
  wire seg_13_19_sp4_v_b_3_50943;
  wire seg_13_19_sp4_v_b_6_50948;
  wire seg_13_19_sp4_v_b_7_50947;
  wire seg_13_19_sp4_v_b_9_50949;
  wire seg_13_1_glb_netwk_0_5;
  wire seg_13_1_glb_netwk_4_9;
  wire seg_13_1_local_g0_3_52784;
  wire seg_13_1_local_g0_4_52785;
  wire seg_13_1_local_g1_2_52791;
  wire seg_13_1_local_g1_3_52792;
  wire seg_13_1_local_g1_4_52793;
  wire seg_13_1_lutff_3_out_48911;
  wire seg_13_1_lutff_5_out_48913;
  wire seg_13_1_neigh_op_top_2_49038;
  wire seg_13_1_neigh_op_top_3_49039;
  wire seg_13_1_neigh_op_top_4_49040;
  wire seg_13_1_sp12_v_b_22_52762;
  wire seg_13_1_sp4_h_r_20_49059;
  wire seg_13_1_sp4_h_r_22_49051;
  wire seg_13_1_sp4_h_r_44_41397;
  wire seg_13_1_sp4_v_b_38_49092;
  wire seg_13_1_sp4_v_b_4_49094;
  wire seg_13_22_sp4_v_b_2_51313;
  wire seg_13_22_sp4_v_b_6_51317;
  wire seg_13_23_sp12_v_b_0_54144;
  wire seg_13_26_sp4_v_b_10_51813;
  wire seg_13_26_sp4_v_b_2_51805;
  wire seg_13_2_glb_netwk_0_5;
  wire seg_13_2_glb_netwk_4_9;
  wire seg_13_2_local_g0_4_52948;
  wire seg_13_2_local_g1_0_52952;
  wire seg_13_2_local_g1_2_52954;
  wire seg_13_2_local_g1_3_52955;
  wire seg_13_2_local_g1_7_52959;
  wire seg_13_2_local_g2_3_52963;
  wire seg_13_2_local_g3_2_52970;
  wire seg_13_2_local_g3_3_52971;
  wire seg_13_2_lutff_0_out_49036;
  wire seg_13_2_lutff_1_out_49037;
  wire seg_13_2_lutff_2_out_49038;
  wire seg_13_2_lutff_3_out_49039;
  wire seg_13_2_lutff_4_out_49040;
  wire seg_13_2_neigh_op_bnl_2_45079;
  wire seg_13_2_neigh_op_bnl_3_45080;
  wire seg_13_2_neigh_op_bot_3_48911;
  wire seg_13_2_neigh_op_top_7_49202;
  wire seg_13_2_sp4_h_l_41_37720;
  wire seg_13_2_sp4_h_l_47_37716;
  wire seg_13_2_sp4_r_v_b_25_52921;
  wire seg_13_2_sp4_r_v_b_37_53051;
  wire seg_13_2_sp4_v_b_10_49076;
  wire seg_13_2_sp4_v_b_6_49071;
  wire seg_13_2_sp4_v_b_8_49074;
  wire seg_13_2_sp4_v_b_9_49073;
  wire seg_13_30_sp4_v_b_10_52305;
  wire seg_13_30_sp4_v_b_1_52294;
  wire seg_13_31_local_g0_3_56527;
  wire seg_13_31_local_g1_0_56532;
  wire seg_13_31_local_g1_0_56532_i1;
  wire seg_13_31_local_g1_0_56532_i2;
  wire seg_13_31_local_g1_0_56532_i3;
  wire seg_13_31_local_g1_1_56533;
  wire seg_13_31_span12_vert_8_55620;
  wire seg_13_31_span4_vert_41_56507;
  wire seg_13_31_span4_vert_43_56509;
  wire seg_13_3_glb_netwk_0_5;
  wire seg_13_3_glb_netwk_4_9;
  wire seg_13_3_local_g0_0_53067;
  wire seg_13_3_local_g0_1_53068;
  wire seg_13_3_local_g0_3_53070;
  wire seg_13_3_local_g0_6_53073;
  wire seg_13_3_local_g0_7_53074;
  wire seg_13_3_local_g1_5_53080;
  wire seg_13_3_local_g2_0_53083;
  wire seg_13_3_local_g2_4_53087;
  wire seg_13_3_local_g2_5_53088;
  wire seg_13_3_local_g3_1_53092;
  wire seg_13_3_local_g3_2_53093;
  wire seg_13_3_lutff_0_out_49195;
  wire seg_13_3_lutff_1_out_49196;
  wire seg_13_3_lutff_2_out_49197;
  wire seg_13_3_lutff_4_out_49199;
  wire seg_13_3_lutff_6_out_49201;
  wire seg_13_3_lutff_7_out_49202;
  wire seg_13_3_neigh_op_tnl_5_45492;
  wire seg_13_3_neigh_op_tnr_2_53151;
  wire seg_13_3_sp4_h_l_37_37837;
  wire seg_13_3_sp4_h_r_10_53163;
  wire seg_13_3_sp4_h_r_16_49337;
  wire seg_13_3_sp4_h_r_1_53162;
  wire seg_13_3_sp4_h_r_2_53165;
  wire seg_13_3_sp4_h_r_8_53171;
  wire seg_13_3_sp4_r_v_b_35_53060;
  wire seg_13_3_sp4_v_b_11_49089;
  wire seg_13_3_sp4_v_b_17_49096;
  wire seg_13_3_sp4_v_b_1_49078;
  wire seg_13_3_sp4_v_b_21_49100;
  wire seg_13_3_sp4_v_b_22_49101;
  wire seg_13_3_sp4_v_b_23_49102;
  wire seg_13_3_sp4_v_b_33_49227;
  wire seg_13_3_sp4_v_b_34_49230;
  wire seg_13_3_sp4_v_t_38_49467;
  wire seg_13_4_glb_netwk_0_5;
  wire seg_13_4_glb_netwk_4_9;
  wire seg_13_4_local_g0_2_53192;
  wire seg_13_4_local_g0_3_53193;
  wire seg_13_4_local_g0_4_53194;
  wire seg_13_4_local_g0_5_53195;
  wire seg_13_4_local_g1_0_53198;
  wire seg_13_4_local_g1_1_53199;
  wire seg_13_4_local_g1_2_53200;
  wire seg_13_4_local_g1_3_53201;
  wire seg_13_4_local_g1_5_53203;
  wire seg_13_4_local_g2_0_53206;
  wire seg_13_4_local_g2_1_53207;
  wire seg_13_4_local_g2_4_53210;
  wire seg_13_4_local_g2_5_53211;
  wire seg_13_4_local_g3_3_53217;
  wire seg_13_4_lutff_0_out_49318;
  wire seg_13_4_lutff_3_out_49321;
  wire seg_13_4_lutff_4_out_49322;
  wire seg_13_4_lutff_5_out_49323;
  wire seg_13_4_lutff_6_out_49324;
  wire seg_13_4_sp12_h_r_10_34126;
  wire seg_13_4_sp4_h_l_40_37967;
  wire seg_13_4_sp4_h_l_41_37966;
  wire seg_13_4_sp4_h_r_11_53287;
  wire seg_13_4_sp4_h_r_16_49460;
  wire seg_13_4_sp4_h_r_20_49464;
  wire seg_13_4_sp4_h_r_22_49456;
  wire seg_13_4_sp4_h_r_28_45628;
  wire seg_13_4_sp4_h_r_32_45632;
  wire seg_13_4_sp4_h_r_36_41792;
  wire seg_13_4_sp4_h_r_38_41796;
  wire seg_13_4_sp4_h_r_3_53289;
  wire seg_13_4_sp4_h_r_4_53290;
  wire seg_13_4_sp4_h_r_5_53291;
  wire seg_13_4_sp4_h_r_8_53294;
  wire seg_13_4_sp4_h_r_9_53295;
  wire seg_13_4_sp4_r_v_b_13_53051;
  wire seg_13_4_sp4_r_v_b_15_53053;
  wire seg_13_4_sp4_r_v_b_1_52921;
  wire seg_13_4_sp4_r_v_b_35_53183;
  wire seg_13_4_sp4_r_v_b_41_53301;
  wire seg_13_4_sp4_v_b_0_49091;
  wire seg_13_4_sp4_v_b_1_49090;
  wire seg_13_4_sp4_v_b_27_49344;
  wire seg_13_4_sp4_v_b_2_49093;
  wire seg_13_4_sp4_v_b_33_49350;
  wire seg_13_4_sp4_v_b_38_49467;
  wire seg_13_4_sp4_v_b_3_49092;
  wire seg_13_4_sp4_v_b_40_49469;
  wire seg_13_4_sp4_v_b_4_49096;
  wire seg_13_4_sp4_v_t_38_49590;
  wire seg_13_5_glb_netwk_0_5;
  wire seg_13_5_local_g0_2_53315;
  wire seg_13_5_local_g1_1_53322;
  wire seg_13_5_local_g1_3_53324;
  wire seg_13_5_local_g2_2_53331;
  wire seg_13_5_local_g2_3_53332;
  wire seg_13_5_lutff_0_out_49441;
  wire seg_13_5_lutff_1_out_49442;
  wire seg_13_5_neigh_op_bot_3_49321;
  wire seg_13_5_sp4_h_l_38_38088;
  wire seg_13_5_sp4_h_l_39_38087;
  wire seg_13_5_sp4_h_r_17_49582;
  wire seg_13_5_sp4_h_r_34_45747;
  wire seg_13_5_sp4_r_v_b_45_53428;
  wire seg_13_5_sp4_v_b_10_49230;
  wire seg_13_5_sp4_v_b_1_49219;
  wire seg_13_5_sp4_v_b_26_49468;
  wire seg_13_5_sp4_v_b_35_49475;
  wire seg_13_5_sp4_v_b_4_49224;
  wire seg_13_6_glb_netwk_0_5;
  wire seg_13_6_glb_netwk_7_12;
  wire seg_13_6_local_g0_3_53439;
  wire seg_13_6_local_g0_5_53441;
  wire seg_13_6_local_g1_1_53445;
  wire seg_13_6_local_g1_6_53450;
  wire seg_13_6_local_g1_7_53451;
  wire seg_13_6_local_g2_1_53453;
  wire seg_13_6_local_g2_2_53454;
  wire seg_13_6_local_g2_3_53455;
  wire seg_13_6_local_g2_6_53458;
  wire seg_13_6_local_g3_2_53462;
  wire seg_13_6_local_g3_7_53467;
  wire seg_13_6_neigh_op_bot_1_49442;
  wire seg_13_6_neigh_op_tnl_1_45857;
  wire seg_13_6_sp4_h_r_0_53530;
  wire seg_13_6_sp4_h_r_10_53532;
  wire seg_13_6_sp4_h_r_15_49703;
  wire seg_13_6_sp4_h_r_20_49710;
  wire seg_13_6_sp4_h_r_26_45872;
  wire seg_13_6_sp4_h_r_27_45873;
  wire seg_13_6_sp4_h_r_2_53534;
  wire seg_13_6_sp4_h_r_30_45876;
  wire seg_13_6_sp4_h_r_44_42048;
  wire seg_13_6_sp4_h_r_4_53536;
  wire seg_13_6_sp4_h_r_8_53540;
  wire seg_13_6_sp4_r_v_b_18_53302;
  wire seg_13_6_sp4_r_v_b_27_53421;
  wire seg_13_6_sp4_r_v_b_7_53179;
  wire seg_13_6_sp4_v_b_0_49343;
  wire seg_13_6_sp4_v_b_21_49474;
  wire seg_13_6_sp4_v_b_22_49475;
  wire seg_13_6_sp4_v_b_30_49595;
  wire seg_13_6_sp4_v_b_39_49714;
  wire seg_13_6_sp4_v_b_5_49346;
  wire seg_13_6_sp4_v_t_38_49836;
  wire seg_13_7_glb_netwk_0_5;
  wire seg_13_7_local_g0_0_53559;
  wire seg_13_7_local_g0_5_53564;
  wire seg_13_7_local_g0_7_53566;
  wire seg_13_7_local_g1_0_53567;
  wire seg_13_7_local_g1_2_53569;
  wire seg_13_7_local_g1_3_53570;
  wire seg_13_7_local_g2_3_53578;
  wire seg_13_7_local_g2_4_53579;
  wire seg_13_7_local_g2_5_53580;
  wire seg_13_7_local_g3_1_53584;
  wire seg_13_7_local_g3_3_53586;
  wire seg_13_7_local_g3_4_53587;
  wire seg_13_7_local_g3_5_53588;
  wire seg_13_7_local_g3_6_53589;
  wire seg_13_7_local_g3_7_53590;
  wire seg_13_7_lutff_0_out_49687;
  wire seg_13_7_lutff_3_out_49690;
  wire seg_13_7_lutff_6_out_49693;
  wire seg_13_7_neigh_op_lft_0_45856;
  wire seg_13_7_neigh_op_lft_7_45863;
  wire seg_13_7_neigh_op_rgt_6_53524;
  wire seg_13_7_sp4_h_l_40_38336;
  wire seg_13_7_sp4_h_r_11_53656;
  wire seg_13_7_sp4_h_r_14_49827;
  wire seg_13_7_sp4_h_r_1_53654;
  wire seg_13_7_sp4_h_r_2_53657;
  wire seg_13_7_sp4_h_r_31_46000;
  wire seg_13_7_sp4_h_r_36_42161;
  wire seg_13_7_sp4_r_v_b_13_53420;
  wire seg_13_7_sp4_r_v_b_17_53424;
  wire seg_13_7_sp4_r_v_b_19_53426;
  wire seg_13_7_sp4_r_v_b_21_53428;
  wire seg_13_7_sp4_r_v_b_37_53666;
  wire seg_13_7_sp4_r_v_b_41_53670;
  wire seg_13_7_sp4_r_v_b_43_53672;
  wire seg_13_7_sp4_v_b_13_49589;
  wire seg_13_7_sp4_v_b_16_49592;
  wire seg_13_7_sp4_v_b_1_49465;
  wire seg_13_7_sp4_v_b_2_49468;
  wire seg_13_7_sp4_v_b_35_49721;
  wire seg_13_7_sp4_v_b_3_49467;
  wire seg_13_7_sp4_v_t_43_49964;
  wire seg_13_8_glb_netwk_0_5;
  wire seg_13_8_glb_netwk_1_6;
  wire seg_13_8_glb_netwk_4_9;
  wire seg_13_8_local_g0_0_53682;
  wire seg_13_8_local_g0_2_53684;
  wire seg_13_8_local_g0_3_53685;
  wire seg_13_8_local_g0_4_53686;
  wire seg_13_8_local_g0_5_53687;
  wire seg_13_8_local_g0_6_53688;
  wire seg_13_8_local_g1_1_53691;
  wire seg_13_8_local_g1_2_53692;
  wire seg_13_8_local_g1_3_53693;
  wire seg_13_8_local_g1_5_53695;
  wire seg_13_8_local_g1_6_53696;
  wire seg_13_8_local_g2_1_53699;
  wire seg_13_8_local_g2_3_53701;
  wire seg_13_8_local_g2_4_53702;
  wire seg_13_8_local_g2_5_53703;
  wire seg_13_8_local_g3_5_53711;
  wire seg_13_8_local_g3_6_53712;
  wire seg_13_8_lutff_5_out_49815;
  wire seg_13_8_lutff_6_out_49816;
  wire seg_13_8_neigh_op_bot_3_49690;
  wire seg_13_8_neigh_op_bot_6_49693;
  wire seg_13_8_neigh_op_top_2_49935;
  wire seg_13_8_neigh_op_top_5_49938;
  wire seg_13_8_sp4_h_l_38_38457;
  wire seg_13_8_sp4_h_l_43_38460;
  wire seg_13_8_sp4_h_r_0_53776;
  wire seg_13_8_sp4_h_r_11_53779;
  wire seg_13_8_sp4_h_r_12_49946;
  wire seg_13_8_sp4_h_r_18_49954;
  wire seg_13_8_sp4_h_r_19_49953;
  wire seg_13_8_sp4_h_r_20_49956;
  wire seg_13_8_sp4_h_r_24_46114;
  wire seg_13_8_sp4_h_r_2_53780;
  wire seg_13_8_sp4_h_r_30_46122;
  wire seg_13_8_sp4_h_r_32_46124;
  wire seg_13_8_sp4_h_r_7_53785;
  wire seg_13_8_sp4_r_v_b_1_53419;
  wire seg_13_8_sp4_r_v_b_35_53675;
  wire seg_13_8_sp4_r_v_b_9_53427;
  wire seg_13_8_sp4_v_b_21_49720;
  wire seg_13_8_sp4_v_b_30_49841;
  wire seg_13_8_sp4_v_b_35_49844;
  wire seg_13_8_sp4_v_b_37_49958;
  wire seg_13_8_sp4_v_b_44_49965;
  wire seg_13_8_sp4_v_b_9_49596;
  wire seg_13_8_sp4_v_t_38_50082;
  wire seg_13_8_sp4_v_t_43_50087;
  wire seg_13_9_glb_netwk_0_5;
  wire seg_13_9_local_g0_6_53811;
  wire seg_13_9_local_g1_3_53816;
  wire seg_13_9_local_g3_3_53832;
  wire seg_13_9_lutff_2_out_49935;
  wire seg_13_9_lutff_5_out_49938;
  wire seg_13_9_sp4_h_l_47_38577;
  wire seg_13_9_sp4_h_r_11_53902;
  wire seg_13_9_sp4_h_r_14_50073;
  wire seg_13_9_sp4_h_r_7_53908;
  wire seg_13_9_sp4_v_b_35_49967;
  wire seg_13_9_sp4_v_t_40_50207;
  wire seg_14_0_span4_horz_r_0_56601;
  wire seg_14_10_glb_netwk_0_5;
  wire seg_14_10_glb_netwk_4_9;
  wire seg_14_10_local_g0_1_57759;
  wire seg_14_10_local_g0_2_57760;
  wire seg_14_10_local_g1_5_57771;
  wire seg_14_10_local_g1_7_57773;
  wire seg_14_10_local_g2_0_57774;
  wire seg_14_10_local_g2_4_57778;
  wire seg_14_10_local_g2_7_57781;
  wire seg_14_10_local_g3_0_57782;
  wire seg_14_10_local_g3_4_57786;
  wire seg_14_10_sp12_h_r_2_54019;
  wire seg_14_10_sp4_h_l_39_42533;
  wire seg_14_10_sp4_h_l_42_42538;
  wire seg_14_10_sp4_h_l_43_42537;
  wire seg_14_10_sp4_h_r_0_57852;
  wire seg_14_10_sp4_h_r_10_57854;
  wire seg_14_10_sp4_h_r_13_54022;
  wire seg_14_10_sp4_h_r_14_54027;
  wire seg_14_10_sp4_h_r_16_54029;
  wire seg_14_10_sp4_h_r_18_54031;
  wire seg_14_10_sp4_h_r_1_57853;
  wire seg_14_10_sp4_h_r_20_54033;
  wire seg_14_10_sp4_h_r_22_54025;
  wire seg_14_10_sp4_h_r_36_46361;
  wire seg_14_10_sp4_h_r_47_46362;
  wire seg_14_10_sp4_h_r_7_57861;
  wire seg_14_10_sp4_h_r_8_57862;
  wire seg_14_10_sp4_h_r_9_57863;
  wire seg_14_10_sp4_r_v_b_13_57619;
  wire seg_14_10_sp4_r_v_b_16_57622;
  wire seg_14_10_sp4_r_v_b_27_57743;
  wire seg_14_10_sp4_r_v_b_29_57745;
  wire seg_14_10_sp4_r_v_b_31_57747;
  wire seg_14_10_sp4_r_v_b_35_57751;
  wire seg_14_10_sp4_v_b_0_53666;
  wire seg_14_10_sp4_v_b_17_53793;
  wire seg_14_10_sp4_v_b_32_53920;
  wire seg_14_10_sp4_v_b_36_54034;
  wire seg_14_10_sp4_v_b_8_53674;
  wire seg_14_10_sp4_v_t_38_54159;
  wire seg_14_10_sp4_v_t_39_54160;
  wire seg_14_11_glb_netwk_0_5;
  wire seg_14_11_local_g0_2_57883;
  wire seg_14_11_local_g0_3_57884;
  wire seg_14_11_local_g1_1_57890;
  wire seg_14_11_local_g1_4_57893;
  wire seg_14_11_local_g1_7_57896;
  wire seg_14_11_sp4_h_l_40_42659;
  wire seg_14_11_sp4_h_r_19_54153;
  wire seg_14_11_sp4_h_r_24_50314;
  wire seg_14_11_sp4_h_r_4_57981;
  wire seg_14_11_sp4_h_r_5_57982;
  wire seg_14_11_sp4_r_v_b_15_57744;
  wire seg_14_11_sp4_r_v_b_17_57746;
  wire seg_14_11_sp4_r_v_b_1_57618;
  wire seg_14_11_sp4_r_v_b_23_57752;
  wire seg_14_11_sp4_v_b_1_53788;
  wire seg_14_11_sp4_v_b_23_53922;
  wire seg_14_11_sp4_v_b_2_53791;
  wire seg_14_11_sp4_v_t_43_54287;
  wire seg_14_12_glb_netwk_0_5;
  wire seg_14_12_glb_netwk_4_9;
  wire seg_14_12_local_g1_0_58012;
  wire seg_14_12_lutff_4_out_54137;
  wire seg_14_12_neigh_op_bnr_0_57840;
  wire seg_14_12_sp4_h_r_11_58101;
  wire seg_14_12_sp4_h_r_6_58106;
  wire seg_14_12_sp4_v_b_11_53921;
  wire seg_14_12_sp4_v_b_1_53911;
  wire seg_14_12_sp4_v_b_40_54284;
  wire seg_14_12_sp4_v_b_8_53920;
  wire seg_14_12_sp4_v_t_42_54409;
  wire seg_14_13_glb_netwk_0_5;
  wire seg_14_13_glb_netwk_4_9;
  wire seg_14_13_local_g0_4_58131;
  wire seg_14_13_local_g0_6_58133;
  wire seg_14_13_local_g1_4_58139;
  wire seg_14_13_local_g2_0_58143;
  wire seg_14_13_local_g2_1_58144;
  wire seg_14_13_local_g2_2_58145;
  wire seg_14_13_local_g2_4_58147;
  wire seg_14_13_local_g3_0_58151;
  wire seg_14_13_local_g3_1_58152;
  wire seg_14_13_local_g3_3_58154;
  wire seg_14_13_local_g3_4_58155;
  wire seg_14_13_lutff_0_out_54256;
  wire seg_14_13_lutff_1_out_54257;
  wire seg_14_13_lutff_3_out_54259;
  wire seg_14_13_lutff_4_out_54260;
  wire seg_14_13_lutff_6_out_54262;
  wire seg_14_13_neigh_op_bot_4_54137;
  wire seg_14_13_neigh_op_tnr_4_58213;
  wire seg_14_13_sp12_h_r_12_35232;
  wire seg_14_13_sp12_v_b_12_57482;
  wire seg_14_13_sp4_h_l_36_42899;
  wire seg_14_13_sp4_h_r_0_58221;
  wire seg_14_13_sp4_h_r_10_58223;
  wire seg_14_13_sp4_h_r_14_54396;
  wire seg_14_13_sp4_h_r_1_58222;
  wire seg_14_13_sp4_h_r_24_50560;
  wire seg_14_13_sp4_h_r_26_50564;
  wire seg_14_13_sp4_h_r_36_46730;
  wire seg_14_13_sp4_h_r_46_46732;
  wire seg_14_13_sp4_h_r_5_58228;
  wire seg_14_13_sp4_r_v_b_21_57996;
  wire seg_14_13_sp4_r_v_b_29_58114;
  wire seg_14_13_sp4_r_v_b_31_58116;
  wire seg_14_13_sp4_r_v_b_33_58118;
  wire seg_14_13_sp4_r_v_b_39_58236;
  wire seg_14_13_sp4_v_b_11_54044;
  wire seg_14_13_sp4_v_b_32_54289;
  wire seg_14_13_sp4_v_b_44_54411;
  wire seg_14_14_glb_netwk_0_5;
  wire seg_14_14_glb_netwk_1_6;
  wire seg_14_14_glb_netwk_4_9;
  wire seg_14_14_local_g0_0_58250;
  wire seg_14_14_local_g0_1_58251;
  wire seg_14_14_local_g0_3_58253;
  wire seg_14_14_local_g0_4_58254;
  wire seg_14_14_local_g1_6_58264;
  wire seg_14_14_local_g2_2_58268;
  wire seg_14_14_local_g2_4_58270;
  wire seg_14_14_local_g2_7_58273;
  wire seg_14_14_local_g3_0_58274;
  wire seg_14_14_local_g3_1_58275;
  wire seg_14_14_lutff_0_out_54379;
  wire seg_14_14_lutff_2_out_54381;
  wire seg_14_14_lutff_4_out_54383;
  wire seg_14_14_lutff_5_out_54384;
  wire seg_14_14_lutff_6_out_54385;
  wire seg_14_14_lutff_7_out_54386;
  wire seg_14_14_neigh_op_bot_3_54259;
  wire seg_14_14_neigh_op_bot_6_54262;
  wire seg_14_14_neigh_op_lft_1_50549;
  wire seg_14_14_sp12_v_b_12_57605;
  wire seg_14_14_sp4_h_l_40_43028;
  wire seg_14_14_sp4_h_r_10_58346;
  wire seg_14_14_sp4_h_r_20_54525;
  wire seg_14_14_sp4_h_r_30_50691;
  wire seg_14_14_sp4_h_r_3_58349;
  wire seg_14_14_sp4_h_r_4_58350;
  wire seg_14_14_sp4_h_r_8_58354;
  wire seg_14_14_sp4_r_v_b_1_57987;
  wire seg_14_14_sp4_r_v_b_33_58241;
  wire seg_14_14_sp4_r_v_b_37_58357;
  wire seg_14_14_sp4_r_v_b_41_58361;
  wire seg_14_14_sp4_r_v_b_43_58363;
  wire seg_14_14_sp4_r_v_b_47_58367;
  wire seg_14_14_sp4_v_b_0_54158;
  wire seg_14_14_sp4_v_b_16_54284;
  wire seg_14_14_sp4_v_b_33_54411;
  wire seg_14_14_sp4_v_b_3_54159;
  wire seg_14_14_sp4_v_t_39_54652;
  wire seg_14_15_glb_netwk_0_5;
  wire seg_14_15_glb_netwk_4_9;
  wire seg_14_15_local_g0_0_58373;
  wire seg_14_15_local_g0_2_58375;
  wire seg_14_15_local_g0_5_58378;
  wire seg_14_15_local_g0_7_58380;
  wire seg_14_15_local_g1_4_58385;
  wire seg_14_15_local_g1_5_58386;
  wire seg_14_15_local_g1_6_58387;
  wire seg_14_15_local_g1_7_58388;
  wire seg_14_15_local_g2_4_58393;
  wire seg_14_15_local_g2_7_58396;
  wire seg_14_15_lutff_0_out_54502;
  wire seg_14_15_lutff_2_out_54504;
  wire seg_14_15_lutff_3_out_54505;
  wire seg_14_15_lutff_4_out_54506;
  wire seg_14_15_lutff_5_out_54507;
  wire seg_14_15_lutff_6_out_54508;
  wire seg_14_15_lutff_7_out_54509;
  wire seg_14_15_neigh_op_bot_0_54379;
  wire seg_14_15_neigh_op_bot_2_54381;
  wire seg_14_15_neigh_op_bot_4_54383;
  wire seg_14_15_neigh_op_bot_5_54384;
  wire seg_14_15_neigh_op_bot_6_54385;
  wire seg_14_15_neigh_op_bot_7_54386;
  wire seg_14_15_sp12_v_b_18_58096;
  wire seg_14_15_sp4_h_l_43_43152;
  wire seg_14_15_sp4_h_r_36_46976;
  wire seg_14_15_sp4_r_v_b_15_58236;
  wire seg_14_15_sp4_r_v_b_5_58114;
  wire seg_14_15_sp4_v_b_10_54291;
  wire seg_14_15_sp4_v_b_15_54406;
  wire seg_14_15_sp4_v_b_7_54286;
  wire seg_14_15_sp4_v_b_8_54289;
  wire seg_14_15_sp4_v_t_39_54775;
  wire seg_14_16_glb_netwk_0_5;
  wire seg_14_16_glb_netwk_4_9;
  wire seg_14_16_local_g0_0_58496;
  wire seg_14_16_local_g0_3_58499;
  wire seg_14_16_local_g0_4_58500;
  wire seg_14_16_local_g0_5_58501;
  wire seg_14_16_local_g0_7_58503;
  wire seg_14_16_local_g1_0_58504;
  wire seg_14_16_local_g1_2_58506;
  wire seg_14_16_local_g1_3_58507;
  wire seg_14_16_local_g1_5_58509;
  wire seg_14_16_local_g1_6_58510;
  wire seg_14_16_local_g1_7_58511;
  wire seg_14_16_local_g2_2_58514;
  wire seg_14_16_local_g2_4_58516;
  wire seg_14_16_local_g3_2_58522;
  wire seg_14_16_local_g3_7_58527;
  wire seg_14_16_neigh_op_bot_0_54502;
  wire seg_14_16_neigh_op_bot_3_54505;
  wire seg_14_16_neigh_op_bot_5_54507;
  wire seg_14_16_neigh_op_bot_6_54508;
  wire seg_14_16_neigh_op_bot_7_54509;
  wire seg_14_16_neigh_op_tnr_2_58580;
  wire seg_14_16_neigh_op_top_7_54755;
  wire seg_14_16_sp4_h_l_38_43272;
  wire seg_14_16_sp4_h_r_10_58592;
  wire seg_14_16_sp4_h_r_14_54765;
  wire seg_14_16_sp4_h_r_20_54771;
  wire seg_14_16_sp4_h_r_24_50929;
  wire seg_14_16_sp4_h_r_31_50938;
  wire seg_14_16_sp4_h_r_4_58596;
  wire seg_14_16_sp4_h_r_8_58600;
  wire seg_14_16_sp4_r_v_b_11_58243;
  wire seg_14_16_sp4_r_v_b_27_58481;
  wire seg_14_16_sp4_r_v_b_29_58483;
  wire seg_14_16_sp4_r_v_b_39_58605;
  wire seg_14_16_sp4_v_b_11_54413;
  wire seg_14_16_sp4_v_b_34_54660;
  wire seg_14_16_sp4_v_b_36_54772;
  wire seg_14_16_sp4_v_b_44_54780;
  wire seg_14_16_sp4_v_b_4_54408;
  wire seg_14_16_sp4_v_t_46_54905;
  wire seg_14_17_glb_netwk_0_5;
  wire seg_14_17_glb_netwk_4_9;
  wire seg_14_17_local_g0_1_58620;
  wire seg_14_17_local_g0_2_58621;
  wire seg_14_17_local_g0_7_58626;
  wire seg_14_17_local_g1_3_58630;
  wire seg_14_17_local_g1_6_58633;
  wire seg_14_17_local_g3_3_58646;
  wire seg_14_17_lutff_2_out_54750;
  wire seg_14_17_lutff_3_out_54751;
  wire seg_14_17_lutff_5_out_54753;
  wire seg_14_17_lutff_6_out_54754;
  wire seg_14_17_lutff_7_out_54755;
  wire seg_14_17_neigh_op_top_1_54872;
  wire seg_14_17_neigh_op_top_7_54878;
  wire seg_14_17_sp4_h_r_0_58713;
  wire seg_14_17_sp4_h_r_11_58716;
  wire seg_14_17_sp4_h_r_14_54888;
  wire seg_14_17_sp4_h_r_2_58717;
  wire seg_14_17_sp4_r_v_b_19_58486;
  wire seg_14_17_sp4_r_v_b_3_58358;
  wire seg_14_17_sp4_v_b_1_54526;
  wire seg_14_17_sp4_v_b_7_54532;
  wire seg_14_18_glb_netwk_0_5;
  wire seg_14_18_glb_netwk_1_6;
  wire seg_14_18_glb_netwk_4_9;
  wire seg_14_18_local_g0_0_58742;
  wire seg_14_18_local_g0_1_58743;
  wire seg_14_18_local_g0_3_58745;
  wire seg_14_18_local_g0_5_58747;
  wire seg_14_18_local_g0_6_58748;
  wire seg_14_18_local_g1_0_58750;
  wire seg_14_18_local_g1_1_58751;
  wire seg_14_18_local_g1_2_58752;
  wire seg_14_18_local_g1_3_58753;
  wire seg_14_18_local_g1_4_58754;
  wire seg_14_18_local_g1_6_58756;
  wire seg_14_18_local_g2_3_58761;
  wire seg_14_18_local_g2_6_58764;
  wire seg_14_18_local_g2_7_58765;
  wire seg_14_18_local_g3_2_58768;
  wire seg_14_18_local_g3_3_58769;
  wire seg_14_18_local_g3_4_58770;
  wire seg_14_18_lutff_0_out_54871;
  wire seg_14_18_lutff_1_out_54872;
  wire seg_14_18_lutff_3_out_54874;
  wire seg_14_18_lutff_5_out_54876;
  wire seg_14_18_lutff_7_out_54878;
  wire seg_14_18_neigh_op_bot_5_54753;
  wire seg_14_18_neigh_op_bot_6_54754;
  wire seg_14_18_neigh_op_lft_1_51041;
  wire seg_14_18_neigh_op_lft_2_51042;
  wire seg_14_18_neigh_op_lft_6_51046;
  wire seg_14_18_sp4_h_l_37_43513;
  wire seg_14_18_sp4_h_l_45_43523;
  wire seg_14_18_sp4_h_r_11_58839;
  wire seg_14_18_sp4_h_r_8_58846;
  wire seg_14_18_sp4_h_r_9_58847;
  wire seg_14_18_sp4_r_v_b_11_58489;
  wire seg_14_18_sp4_r_v_b_13_58603;
  wire seg_14_18_sp4_r_v_b_14_58604;
  wire seg_14_18_sp4_r_v_b_15_58605;
  wire seg_14_18_sp4_r_v_b_20_58610;
  wire seg_14_18_sp4_r_v_b_35_58735;
  wire seg_14_18_sp4_r_v_b_3_58481;
  wire seg_14_18_sp4_r_v_b_5_58483;
  wire seg_14_18_sp4_v_b_0_54650;
  wire seg_14_18_sp4_v_b_10_54660;
  wire seg_14_18_sp4_v_b_12_54772;
  wire seg_14_18_sp4_v_b_20_54780;
  wire seg_14_18_sp4_v_b_26_54898;
  wire seg_14_18_sp4_v_b_2_54652;
  wire seg_14_18_sp4_v_b_3_54651;
  wire seg_14_19_glb_netwk_0_5;
  wire seg_14_19_glb_netwk_4_9;
  wire seg_14_19_local_g2_2_58883;
  wire seg_14_19_local_g2_3_58884;
  wire seg_14_19_local_g3_0_58889;
  wire seg_14_19_local_g3_3_58892;
  wire seg_14_19_local_g3_7_58896;
  wire seg_14_19_lutff_3_out_54997;
  wire seg_14_19_sp12_v_b_0_57482;
  wire seg_14_19_sp12_v_b_10_58096;
  wire seg_14_19_sp12_v_b_3_57605;
  wire seg_14_19_sp4_r_v_b_23_58736;
  wire seg_14_19_sp4_v_b_22_54905;
  wire seg_14_1_local_g0_3_56614;
  wire seg_14_1_local_g2_0_56627;
  wire seg_14_1_neigh_op_lft_3_48911;
  wire seg_14_1_neigh_op_tnl_0_49036;
  wire seg_14_1_sp4_h_r_44_45228;
  wire seg_14_1_sp4_v_b_1_52892;
  wire seg_14_2_glb_netwk_0_5;
  wire seg_14_2_glb_netwk_3_8;
  wire seg_14_2_glb_netwk_4_9;
  wire seg_14_2_local_g0_0_56774;
  wire seg_14_2_local_g0_2_56776;
  wire seg_14_2_local_g0_5_56779;
  wire seg_14_2_local_g1_1_56783;
  wire seg_14_2_local_g1_3_56785;
  wire seg_14_2_local_g1_6_56788;
  wire seg_14_2_lutff_0_out_52867;
  wire seg_14_2_lutff_2_out_52869;
  wire seg_14_2_lutff_6_out_52873;
  wire seg_14_2_sp4_h_r_17_53044;
  wire seg_14_2_sp4_h_r_19_53046;
  wire seg_14_2_sp4_h_r_21_53048;
  wire seg_14_2_sp4_r_v_b_39_56883;
  wire seg_14_2_sp4_v_t_46_53183;
  wire seg_14_3_glb_netwk_0_5;
  wire seg_14_3_glb_netwk_3_8;
  wire seg_14_3_glb_netwk_4_9;
  wire seg_14_3_local_g0_3_56900;
  wire seg_14_3_local_g1_2_56907;
  wire seg_14_3_lutff_6_out_53032;
  wire seg_14_3_lutff_7_out_53033;
  wire seg_14_3_sp4_h_l_41_41674;
  wire seg_14_3_sp4_h_r_11_56994;
  wire seg_14_3_sp4_h_r_18_53170;
  wire seg_14_3_sp4_v_t_46_53306;
  wire seg_14_4_glb_netwk_0_5;
  wire seg_14_4_glb_netwk_3_8;
  wire seg_14_4_local_g0_0_57020;
  wire seg_14_4_local_g0_6_57026;
  wire seg_14_4_local_g1_4_57032;
  wire seg_14_4_local_g1_7_57035;
  wire seg_14_4_local_g2_4_57040;
  wire seg_14_4_local_g2_7_57043;
  wire seg_14_4_local_g3_1_57045;
  wire seg_14_4_local_g3_4_57048;
  wire seg_14_4_local_g3_7_57051;
  wire seg_14_4_lutff_0_out_53149;
  wire seg_14_4_lutff_2_out_53151;
  wire seg_14_4_lutff_3_out_53152;
  wire seg_14_4_lutff_5_out_53154;
  wire seg_14_4_neigh_op_bnl_1_49196;
  wire seg_14_4_neigh_op_bot_6_53032;
  wire seg_14_4_neigh_op_bot_7_53033;
  wire seg_14_4_neigh_op_lft_0_49318;
  wire seg_14_4_sp4_h_r_12_53285;
  wire seg_14_4_sp4_h_r_20_53295;
  wire seg_14_4_sp4_h_r_28_49459;
  wire seg_14_4_sp4_h_r_30_49461;
  wire seg_14_4_sp4_h_r_36_45623;
  wire seg_14_4_sp4_h_r_44_45633;
  wire seg_14_4_sp4_r_v_b_15_56883;
  wire seg_14_4_sp4_r_v_b_21_56889;
  wire seg_14_4_sp4_r_v_b_23_56891;
  wire seg_14_4_sp4_r_v_b_25_57003;
  wire seg_14_4_sp4_r_v_b_45_57135;
  wire seg_14_4_sp4_v_b_36_53296;
  wire seg_14_5_glb_netwk_0_5;
  wire seg_14_5_local_g0_0_57143;
  wire seg_14_5_local_g0_2_57145;
  wire seg_14_5_local_g0_3_57146;
  wire seg_14_5_local_g1_1_57152;
  wire seg_14_5_local_g1_4_57155;
  wire seg_14_5_local_g1_5_57156;
  wire seg_14_5_local_g2_0_57159;
  wire seg_14_5_local_g2_1_57160;
  wire seg_14_5_local_g2_3_57162;
  wire seg_14_5_local_g2_4_57163;
  wire seg_14_5_local_g2_6_57165;
  wire seg_14_5_local_g2_7_57166;
  wire seg_14_5_local_g3_1_57168;
  wire seg_14_5_local_g3_3_57170;
  wire seg_14_5_local_g3_5_57172;
  wire seg_14_5_local_g3_6_57173;
  wire seg_14_5_local_g3_7_57174;
  wire seg_14_5_lutff_1_out_53273;
  wire seg_14_5_lutff_2_out_53274;
  wire seg_14_5_lutff_3_out_53275;
  wire seg_14_5_lutff_4_out_53276;
  wire seg_14_5_lutff_5_out_53277;
  wire seg_14_5_lutff_6_out_53278;
  wire seg_14_5_lutff_7_out_53279;
  wire seg_14_5_neigh_op_bnl_3_49321;
  wire seg_14_5_neigh_op_bnl_4_49322;
  wire seg_14_5_neigh_op_bot_0_53149;
  wire seg_14_5_neigh_op_bot_3_53152;
  wire seg_14_5_neigh_op_bot_5_53154;
  wire seg_14_5_sp4_h_r_17_53413;
  wire seg_14_5_sp4_h_r_32_49586;
  wire seg_14_5_sp4_h_r_41_45751;
  wire seg_14_5_sp4_r_v_b_17_57008;
  wire seg_14_5_sp4_v_b_11_53060;
  wire seg_14_5_sp4_v_b_12_53173;
  wire seg_14_5_sp4_v_b_2_53053;
  wire seg_14_5_sp4_v_b_30_53303;
  wire seg_14_5_sp4_v_b_31_53302;
  wire seg_14_5_sp4_v_b_37_53420;
  wire seg_14_5_sp4_v_b_43_53426;
  wire seg_14_6_glb_netwk_0_5;
  wire seg_14_6_glb_netwk_4_9;
  wire seg_14_6_local_g0_0_57266;
  wire seg_14_6_local_g0_3_57269;
  wire seg_14_6_local_g0_4_57270;
  wire seg_14_6_local_g0_7_57273;
  wire seg_14_6_local_g1_1_57275;
  wire seg_14_6_local_g1_2_57276;
  wire seg_14_6_local_g1_3_57277;
  wire seg_14_6_local_g1_4_57278;
  wire seg_14_6_local_g1_5_57279;
  wire seg_14_6_local_g2_0_57282;
  wire seg_14_6_local_g2_6_57288;
  wire seg_14_6_local_g3_0_57290;
  wire seg_14_6_local_g3_4_57294;
  wire seg_14_6_local_g3_5_57295;
  wire seg_14_6_local_g3_6_57296;
  wire seg_14_6_lutff_0_out_53395;
  wire seg_14_6_lutff_3_out_53398;
  wire seg_14_6_lutff_5_out_53400;
  wire seg_14_6_lutff_7_out_53402;
  wire seg_14_6_neigh_op_bnl_0_49441;
  wire seg_14_6_neigh_op_bot_3_53275;
  wire seg_14_6_neigh_op_bot_7_53279;
  wire seg_14_6_neigh_op_rgt_0_57225;
  wire seg_14_6_neigh_op_rgt_4_57229;
  wire seg_14_6_sp12_h_r_0_57356;
  wire seg_14_6_sp4_h_l_39_42041;
  wire seg_14_6_sp4_h_l_42_42046;
  wire seg_14_6_sp4_h_l_44_42048;
  wire seg_14_6_sp4_h_r_0_57360;
  wire seg_14_6_sp4_h_r_2_57364;
  wire seg_14_6_sp4_h_r_44_45879;
  wire seg_14_6_sp4_h_r_4_57366;
  wire seg_14_6_sp4_h_r_8_57370;
  wire seg_14_6_sp4_r_v_b_1_57003;
  wire seg_14_6_sp4_r_v_b_21_57135;
  wire seg_14_6_sp4_v_b_12_53296;
  wire seg_14_6_sp4_v_b_13_53297;
  wire seg_14_6_sp4_v_b_18_53302;
  wire seg_14_6_sp4_v_b_19_53303;
  wire seg_14_6_sp4_v_b_20_53304;
  wire seg_14_6_sp4_v_b_30_53426;
  wire seg_14_6_sp4_v_b_7_53179;
  wire seg_14_7_glb_netwk_0_5;
  wire seg_14_7_glb_netwk_4_9;
  wire seg_14_7_local_g0_7_57396;
  wire seg_14_7_local_g1_5_57402;
  wire seg_14_7_local_g1_7_57404;
  wire seg_14_7_local_g2_2_57407;
  wire seg_14_7_local_g3_3_57416;
  wire seg_14_7_lutff_1_out_53519;
  wire seg_14_7_lutff_5_out_53523;
  wire seg_14_7_lutff_6_out_53524;
  wire seg_14_7_lutff_7_out_53525;
  wire seg_14_7_neigh_op_bot_5_53400;
  wire seg_14_7_neigh_op_rgt_2_57350;
  wire seg_14_7_neigh_op_rgt_3_57351;
  wire seg_14_7_sp4_h_l_36_42161;
  wire seg_14_7_sp4_h_l_37_42160;
  wire seg_14_7_sp4_h_l_38_42165;
  wire seg_14_7_sp4_h_l_43_42168;
  wire seg_14_7_sp4_h_r_11_57486;
  wire seg_14_7_sp4_h_r_12_53654;
  wire seg_14_7_sp4_h_r_23_53655;
  wire seg_14_7_sp4_h_r_28_49828;
  wire seg_14_7_sp4_h_r_38_45996;
  wire seg_14_7_sp4_h_r_5_57490;
  wire seg_14_7_sp4_v_b_1_53296;
  wire seg_14_7_sp4_v_b_44_53673;
  wire seg_14_7_sp4_v_b_4_53301;
  wire seg_14_8_glb_netwk_0_5;
  wire seg_14_8_glb_netwk_4_9;
  wire seg_14_8_local_g0_0_57512;
  wire seg_14_8_local_g0_1_57513;
  wire seg_14_8_local_g0_5_57517;
  wire seg_14_8_local_g1_1_57521;
  wire seg_14_8_local_g1_3_57523;
  wire seg_14_8_local_g1_4_57524;
  wire seg_14_8_local_g1_5_57525;
  wire seg_14_8_local_g2_0_57528;
  wire seg_14_8_local_g3_0_57536;
  wire seg_14_8_local_g3_2_57538;
  wire seg_14_8_local_g3_5_57541;
  wire seg_14_8_lutff_5_out_53646;
  wire seg_14_8_neigh_op_bnl_0_49687;
  wire seg_14_8_neigh_op_bnr_4_57352;
  wire seg_14_8_neigh_op_bot_1_53519;
  wire seg_14_8_neigh_op_bot_5_53523;
  wire seg_14_8_neigh_op_top_0_53764;
  wire seg_14_8_sp4_h_l_37_42283;
  wire seg_14_8_sp4_h_l_44_42294;
  wire seg_14_8_sp4_h_r_0_57606;
  wire seg_14_8_sp4_h_r_10_57608;
  wire seg_14_8_sp4_h_r_11_57609;
  wire seg_14_8_sp4_h_r_12_53777;
  wire seg_14_8_sp4_h_r_17_53782;
  wire seg_14_8_sp4_h_r_1_57607;
  wire seg_14_8_sp4_h_r_21_53786;
  wire seg_14_8_sp4_h_r_22_53779;
  wire seg_14_8_sp4_h_r_2_57610;
  wire seg_14_8_sp4_h_r_38_46119;
  wire seg_14_8_sp4_h_r_40_46121;
  wire seg_14_8_sp4_h_r_46_46117;
  wire seg_14_8_sp4_h_r_5_57613;
  wire seg_14_8_sp4_h_r_8_57616;
  wire seg_14_8_sp4_h_r_9_57617;
  wire seg_14_8_sp4_r_v_b_27_57497;
  wire seg_14_8_sp4_r_v_b_39_57621;
  wire seg_14_8_sp4_r_v_b_47_57629;
  wire seg_14_8_sp4_v_b_20_53550;
  wire seg_14_8_sp4_v_b_22_53552;
  wire seg_14_8_sp4_v_b_29_53669;
  wire seg_14_8_sp4_v_b_32_53674;
  wire seg_14_8_sp4_v_b_34_53676;
  wire seg_14_8_sp4_v_b_36_53788;
  wire seg_14_8_sp4_v_b_46_53798;
  wire seg_14_8_sp4_v_t_42_53917;
  wire seg_14_9_glb_netwk_0_5;
  wire seg_14_9_local_g0_0_57635;
  wire seg_14_9_local_g0_1_57636;
  wire seg_14_9_local_g0_2_57637;
  wire seg_14_9_local_g0_4_57639;
  wire seg_14_9_local_g1_0_57643;
  wire seg_14_9_local_g1_1_57644;
  wire seg_14_9_local_g1_3_57646;
  wire seg_14_9_lutff_0_out_53764;
  wire seg_14_9_lutff_1_out_53765;
  wire seg_14_9_neigh_op_bnr_2_57473;
  wire seg_14_9_neigh_op_bnr_4_57475;
  wire seg_14_9_sp4_h_l_41_42412;
  wire seg_14_9_sp4_h_l_45_42416;
  wire seg_14_9_sp4_h_r_0_57729;
  wire seg_14_9_sp4_h_r_10_57731;
  wire seg_14_9_sp4_h_r_16_53906;
  wire seg_14_9_sp4_h_r_3_57734;
  wire seg_14_9_sp4_h_r_9_57740;
  wire seg_14_9_sp4_r_v_b_27_57620;
  wire seg_14_9_sp4_r_v_b_45_57750;
  wire seg_14_9_sp4_v_b_11_53552;
  wire seg_14_9_sp4_v_b_16_53669;
  wire seg_14_9_sp4_v_b_17_53670;
  wire seg_14_9_sp4_v_b_9_53550;
  wire seg_15_0_span4_horz_r_0_60431;
  wire seg_15_0_span4_vert_24_56738;
  wire seg_15_10_glb_netwk_0_5;
  wire seg_15_10_glb_netwk_4_9;
  wire seg_15_10_local_g0_0_61588;
  wire seg_15_10_local_g0_6_61594;
  wire seg_15_10_local_g1_0_61596;
  wire seg_15_10_local_g1_1_61597;
  wire seg_15_10_local_g1_6_61602;
  wire seg_15_10_local_g2_2_61606;
  wire seg_15_10_local_g2_3_61607;
  wire seg_15_10_local_g2_6_61610;
  wire seg_15_10_local_g3_2_61614;
  wire seg_15_10_lutff_1_out_57718;
  wire seg_15_10_lutff_2_out_57719;
  wire seg_15_10_lutff_3_out_57720;
  wire seg_15_10_lutff_6_out_57723;
  wire seg_15_10_neigh_op_top_0_57840;
  wire seg_15_10_sp4_h_r_0_61682;
  wire seg_15_10_sp4_h_r_14_57857;
  wire seg_15_10_sp4_h_r_26_54026;
  wire seg_15_10_sp4_h_r_2_61686;
  wire seg_15_10_sp4_h_r_30_54030;
  wire seg_15_10_sp4_v_b_11_57505;
  wire seg_15_10_sp4_v_b_8_57504;
  wire seg_15_10_sp4_v_t_39_57990;
  wire seg_15_11_glb_netwk_0_5;
  wire seg_15_11_glb_netwk_4_9;
  wire seg_15_11_local_g0_2_61713;
  wire seg_15_11_local_g0_3_61714;
  wire seg_15_11_local_g1_1_61720;
  wire seg_15_11_local_g1_4_61723;
  wire seg_15_11_local_g1_5_61724;
  wire seg_15_11_local_g1_6_61725;
  wire seg_15_11_local_g2_4_61731;
  wire seg_15_11_local_g2_6_61733;
  wire seg_15_11_local_g2_7_61734;
  wire seg_15_11_local_g3_1_61736;
  wire seg_15_11_local_g3_2_61737;
  wire seg_15_11_local_g3_7_61742;
  wire seg_15_11_lutff_0_out_57840;
  wire seg_15_11_lutff_1_out_57841;
  wire seg_15_11_lutff_2_out_57842;
  wire seg_15_11_lutff_3_out_57843;
  wire seg_15_11_lutff_4_out_57844;
  wire seg_15_11_lutff_7_out_57847;
  wire seg_15_11_neigh_op_bot_1_57718;
  wire seg_15_11_neigh_op_bot_2_57719;
  wire seg_15_11_neigh_op_bot_3_57720;
  wire seg_15_11_neigh_op_bot_6_57723;
  wire seg_15_11_neigh_op_rgt_6_61676;
  wire seg_15_11_neigh_op_rgt_7_61677;
  wire seg_15_11_sp4_h_l_46_46486;
  wire seg_15_11_sp4_h_r_0_61805;
  wire seg_15_11_sp4_h_r_16_57982;
  wire seg_15_11_sp4_h_r_22_57978;
  wire seg_15_11_sp4_h_r_28_54151;
  wire seg_15_11_sp4_h_r_31_54154;
  wire seg_15_11_sp4_h_r_42_50323;
  wire seg_15_11_sp4_h_r_5_61812;
  wire seg_15_11_sp4_r_v_b_33_61702;
  wire seg_15_11_sp4_r_v_b_45_61826;
  wire seg_15_11_sp4_r_v_b_5_61452;
  wire seg_15_11_sp4_v_b_0_57619;
  wire seg_15_11_sp4_v_b_10_57629;
  wire seg_15_11_sp4_v_b_12_57741;
  wire seg_15_11_sp4_v_b_20_57749;
  wire seg_15_11_sp4_v_b_2_57621;
  wire seg_15_11_sp4_v_b_44_57995;
  wire seg_15_11_sp4_v_b_7_57624;
  wire seg_15_11_sp4_v_b_9_57626;
  wire seg_15_11_sp4_v_t_38_58112;
  wire seg_15_11_sp4_v_t_41_58115;
  wire seg_15_11_sp4_v_t_46_58120;
  wire seg_15_12_glb_netwk_0_5;
  wire seg_15_12_glb_netwk_4_9;
  wire seg_15_12_local_g0_7_61841;
  wire seg_15_12_local_g1_1_61843;
  wire seg_15_12_local_g1_7_61849;
  wire seg_15_12_local_g2_1_61851;
  wire seg_15_12_local_g2_2_61852;
  wire seg_15_12_local_g2_4_61854;
  wire seg_15_12_local_g2_7_61857;
  wire seg_15_12_local_g3_6_61864;
  wire seg_15_12_local_g3_7_61865;
  wire seg_15_12_lutff_1_out_57964;
  wire seg_15_12_lutff_2_out_57965;
  wire seg_15_12_lutff_3_out_57966;
  wire seg_15_12_lutff_4_out_57967;
  wire seg_15_12_lutff_6_out_57969;
  wire seg_15_12_lutff_7_out_57970;
  wire seg_15_12_neigh_op_bot_7_57847;
  wire seg_15_12_neigh_op_top_7_58093;
  wire seg_15_12_sp4_h_r_9_61939;
  wire seg_15_12_sp4_r_v_b_33_61825;
  wire seg_15_12_sp4_r_v_b_47_61951;
  wire seg_15_12_sp4_v_b_10_57752;
  wire seg_15_12_sp4_v_b_11_57751;
  wire seg_15_12_sp4_v_b_1_57741;
  wire seg_15_12_sp4_v_b_25_57987;
  wire seg_15_12_sp4_v_b_26_57990;
  wire seg_15_12_sp4_v_b_2_57744;
  wire seg_15_12_sp4_v_b_30_57994;
  wire seg_15_12_sp4_v_b_34_57998;
  wire seg_15_12_sp4_v_b_36_58110;
  wire seg_15_12_sp4_v_b_3_57743;
  wire seg_15_12_sp4_v_b_4_57746;
  wire seg_15_12_sp4_v_b_5_57745;
  wire seg_15_12_sp4_v_b_7_57747;
  wire seg_15_12_sp4_v_b_8_57750;
  wire seg_15_12_sp4_v_t_36_58233;
  wire seg_15_13_glb_netwk_0_5;
  wire seg_15_13_glb_netwk_4_9;
  wire seg_15_13_local_g0_5_61962;
  wire seg_15_13_local_g1_3_61968;
  wire seg_15_13_local_g2_2_61975;
  wire seg_15_13_local_g2_3_61976;
  wire seg_15_13_local_g3_1_61982;
  wire seg_15_13_local_g3_4_61985;
  wire seg_15_13_local_g3_5_61986;
  wire seg_15_13_local_g3_6_61987;
  wire seg_15_13_lutff_1_out_58087;
  wire seg_15_13_lutff_2_out_58088;
  wire seg_15_13_lutff_3_out_58089;
  wire seg_15_13_lutff_5_out_58091;
  wire seg_15_13_lutff_7_out_58093;
  wire seg_15_13_neigh_op_rgt_1_61917;
  wire seg_15_13_neigh_op_rgt_2_61918;
  wire seg_15_13_neigh_op_rgt_3_61919;
  wire seg_15_13_neigh_op_rgt_4_61920;
  wire seg_15_13_neigh_op_rgt_5_61921;
  wire seg_15_13_neigh_op_rgt_6_61922;
  wire seg_15_13_neigh_op_top_5_58214;
  wire seg_15_13_sp4_h_r_40_50567;
  wire seg_15_13_sp4_v_b_19_57994;
  wire seg_15_13_sp4_v_b_28_58115;
  wire seg_15_13_sp4_v_b_2_57867;
  wire seg_15_13_sp4_v_t_38_58358;
  wire seg_15_14_glb_netwk_0_5;
  wire seg_15_14_glb_netwk_4_9;
  wire seg_15_14_local_g0_1_62081;
  wire seg_15_14_local_g0_2_62082;
  wire seg_15_14_local_g0_3_62083;
  wire seg_15_14_local_g0_5_62085;
  wire seg_15_14_local_g1_2_62090;
  wire seg_15_14_local_g1_3_62091;
  wire seg_15_14_local_g1_4_62092;
  wire seg_15_14_local_g1_5_62093;
  wire seg_15_14_local_g2_0_62096;
  wire seg_15_14_local_g2_1_62097;
  wire seg_15_14_local_g3_3_62107;
  wire seg_15_14_local_g3_5_62109;
  wire seg_15_14_lutff_1_out_58210;
  wire seg_15_14_lutff_4_out_58213;
  wire seg_15_14_lutff_5_out_58214;
  wire seg_15_14_neigh_op_bnl_0_54256;
  wire seg_15_14_neigh_op_bot_1_58087;
  wire seg_15_14_neigh_op_bot_2_58088;
  wire seg_15_14_neigh_op_bot_3_58089;
  wire seg_15_14_neigh_op_bot_5_58091;
  wire seg_15_14_neigh_op_tnr_5_62167;
  wire seg_15_14_neigh_op_top_4_58336;
  wire seg_15_14_sp4_h_r_0_62174;
  wire seg_15_14_sp4_h_r_20_58355;
  wire seg_15_14_sp4_h_r_24_54514;
  wire seg_15_14_sp4_h_r_28_54520;
  wire seg_15_14_sp4_h_r_34_54516;
  wire seg_15_14_sp4_h_r_46_50686;
  wire seg_15_14_sp4_h_r_4_62180;
  wire seg_15_14_sp4_r_v_b_19_61947;
  wire seg_15_14_sp4_r_v_b_23_61951;
  wire seg_15_14_sp4_r_v_b_2_61820;
  wire seg_15_14_sp4_r_v_b_3_61819;
  wire seg_15_14_sp4_r_v_b_47_62197;
  wire seg_15_14_sp4_r_v_b_7_61823;
  wire seg_15_14_sp4_r_v_b_9_61825;
  wire seg_15_14_sp4_v_b_10_57998;
  wire seg_15_14_sp4_v_b_11_57997;
  wire seg_15_14_sp4_v_b_12_58110;
  wire seg_15_14_sp4_v_b_13_58111;
  wire seg_15_14_sp4_v_b_4_57992;
  wire seg_15_14_sp4_v_b_8_57996;
  wire seg_15_14_sp4_v_b_9_57995;
  wire seg_15_14_sp4_v_t_43_58486;
  wire seg_15_15_glb_netwk_0_5;
  wire seg_15_15_glb_netwk_4_9;
  wire seg_15_15_local_g1_1_62212;
  wire seg_15_15_local_g1_2_62213;
  wire seg_15_15_local_g1_3_62214;
  wire seg_15_15_local_g3_1_62228;
  wire seg_15_15_local_g3_5_62232;
  wire seg_15_15_local_g3_6_62233;
  wire seg_15_15_lutff_1_out_58333;
  wire seg_15_15_lutff_2_out_58334;
  wire seg_15_15_lutff_3_out_58335;
  wire seg_15_15_lutff_4_out_58336;
  wire seg_15_15_neigh_op_bot_1_58210;
  wire seg_15_15_neigh_op_rgt_6_62168;
  wire seg_15_15_sp4_h_l_44_46986;
  wire seg_15_15_sp4_h_l_46_46978;
  wire seg_15_15_sp4_r_v_b_15_62066;
  wire seg_15_15_sp4_r_v_b_17_62068;
  wire seg_15_15_sp4_r_v_b_3_61942;
  wire seg_15_15_sp4_r_v_b_9_61948;
  wire seg_15_15_sp4_v_b_12_58233;
  wire seg_15_15_sp4_v_b_32_58365;
  wire seg_15_15_sp4_v_b_45_58488;
  wire seg_15_15_sp4_v_b_7_58116;
  wire seg_15_16_glb_netwk_0_5;
  wire seg_15_16_glb_netwk_4_9;
  wire seg_15_16_local_g0_0_62326;
  wire seg_15_16_local_g0_1_62327;
  wire seg_15_16_local_g0_5_62331;
  wire seg_15_16_local_g0_7_62333;
  wire seg_15_16_local_g1_1_62335;
  wire seg_15_16_local_g1_3_62337;
  wire seg_15_16_local_g2_0_62342;
  wire seg_15_16_local_g2_3_62345;
  wire seg_15_16_local_g2_5_62347;
  wire seg_15_16_local_g2_6_62348;
  wire seg_15_16_local_g3_1_62351;
  wire seg_15_16_local_g3_2_62352;
  wire seg_15_16_local_g3_3_62353;
  wire seg_15_16_local_g3_5_62355;
  wire seg_15_16_local_g3_6_62356;
  wire seg_15_16_lutff_1_out_58456;
  wire seg_15_16_lutff_2_out_58457;
  wire seg_15_16_lutff_4_out_58459;
  wire seg_15_16_lutff_5_out_58460;
  wire seg_15_16_lutff_7_out_58462;
  wire seg_15_16_neigh_op_rgt_0_62285;
  wire seg_15_16_neigh_op_rgt_1_62286;
  wire seg_15_16_neigh_op_rgt_6_62291;
  wire seg_15_16_neigh_op_tnr_2_62410;
  wire seg_15_16_sp4_r_v_b_14_62188;
  wire seg_15_16_sp4_v_b_11_58243;
  wire seg_15_16_sp4_v_b_13_58357;
  wire seg_15_16_sp4_v_b_16_58360;
  wire seg_15_16_sp4_v_b_17_58361;
  wire seg_15_16_sp4_v_b_19_58363;
  wire seg_15_16_sp4_v_b_23_58367;
  wire seg_15_16_sp4_v_b_27_58481;
  wire seg_15_16_sp4_v_b_29_58483;
  wire seg_15_16_sp4_v_b_2_58236;
  wire seg_15_16_sp4_v_b_35_58489;
  wire seg_15_16_sp4_v_b_37_58603;
  wire seg_15_16_sp4_v_b_38_58604;
  wire seg_15_16_sp4_v_b_3_58235;
  wire seg_15_16_sp4_v_b_44_58610;
  wire seg_15_16_sp4_v_b_9_58241;
  wire seg_15_17_glb_netwk_0_5;
  wire seg_15_17_glb_netwk_4_9;
  wire seg_15_17_local_g0_0_62449;
  wire seg_15_17_local_g2_1_62466;
  wire seg_15_17_local_g2_2_62467;
  wire seg_15_17_local_g2_3_62468;
  wire seg_15_17_local_g2_5_62470;
  wire seg_15_17_local_g3_7_62480;
  wire seg_15_17_lutff_0_out_58578;
  wire seg_15_17_lutff_2_out_58580;
  wire seg_15_17_lutff_4_out_58582;
  wire seg_15_17_neigh_op_rgt_3_62411;
  wire seg_15_17_neigh_op_tnl_1_54872;
  wire seg_15_17_neigh_op_tnl_5_54876;
  wire seg_15_17_neigh_op_tnl_7_54878;
  wire seg_15_17_sp4_h_r_0_62543;
  wire seg_15_17_sp4_h_r_16_58720;
  wire seg_15_17_sp4_h_r_2_62547;
  wire seg_15_17_sp4_v_b_6_58363;
  wire seg_15_17_sp4_v_b_8_58365;
  wire seg_15_18_glb_netwk_0_5;
  wire seg_15_18_glb_netwk_4_9;
  wire seg_15_18_local_g0_3_62575;
  wire seg_15_18_local_g1_2_62582;
  wire seg_15_18_local_g1_3_62583;
  wire seg_15_18_local_g2_4_62592;
  wire seg_15_18_local_g3_1_62597;
  wire seg_15_18_sp4_h_r_19_58844;
  wire seg_15_18_sp4_r_v_b_12_62432;
  wire seg_15_18_sp4_r_v_b_17_62437;
  wire seg_15_18_sp4_r_v_b_3_62311;
  wire seg_15_18_sp4_v_b_2_58482;
  wire seg_15_18_sp4_v_b_8_58488;
  wire seg_15_1_sp4_h_l_44_45228;
  wire seg_15_1_sp4_h_r_5_60546;
  wire seg_15_2_glb_netwk_0_5;
  wire seg_15_2_glb_netwk_7_12;
  wire seg_15_2_local_g2_7_60627;
  wire seg_15_2_sp4_h_l_47_45378;
  wire seg_15_2_sp4_h_r_11_60701;
  wire seg_15_2_sp4_h_r_1_60699;
  wire seg_15_2_sp4_h_r_39_49211;
  wire seg_15_2_sp4_h_r_5_60705;
  wire seg_15_2_sp4_h_r_8_60708;
  wire seg_15_2_sp4_v_b_28_56757;
  wire seg_15_3_glb_netwk_0_5;
  wire seg_15_3_glb_netwk_4_9;
  wire seg_15_3_local_g0_2_60729;
  wire seg_15_3_local_g0_4_60731;
  wire seg_15_3_lutff_2_out_56858;
  wire seg_15_3_neigh_op_top_2_56981;
  wire seg_15_3_sp4_h_r_12_56992;
  wire seg_15_3_sp4_h_r_40_49337;
  wire seg_15_3_sp4_v_b_0_56738;
  wire seg_15_3_sp4_v_b_1_56739;
  wire seg_15_4_glb_netwk_0_5;
  wire seg_15_4_glb_netwk_4_9;
  wire seg_15_4_local_g0_0_60850;
  wire seg_15_4_local_g0_2_60852;
  wire seg_15_4_local_g1_2_60860;
  wire seg_15_4_local_g2_0_60866;
  wire seg_15_4_local_g2_4_60870;
  wire seg_15_4_local_g3_0_60874;
  wire seg_15_4_local_g3_2_60876;
  wire seg_15_4_local_g3_4_60878;
  wire seg_15_4_local_g3_6_60880;
  wire seg_15_4_lutff_0_out_56979;
  wire seg_15_4_lutff_2_out_56981;
  wire seg_15_4_lutff_7_out_56986;
  wire seg_15_4_neigh_op_lft_2_53151;
  wire seg_15_4_sp4_h_r_24_53284;
  wire seg_15_4_sp4_h_r_26_53288;
  wire seg_15_4_sp4_h_r_28_53290;
  wire seg_15_4_sp4_h_r_30_53292;
  wire seg_15_4_sp4_h_r_32_53294;
  wire seg_15_4_sp4_h_r_34_53286;
  wire seg_15_4_sp4_h_r_40_49460;
  wire seg_15_4_sp4_h_r_42_49462;
  wire seg_15_4_sp4_h_r_6_60952;
  wire seg_15_4_sp4_r_v_b_26_60836;
  wire seg_15_4_sp4_r_v_b_29_60837;
  wire seg_15_4_sp4_r_v_b_39_60959;
  wire seg_15_4_sp4_r_v_b_41_60961;
  wire seg_15_4_sp4_v_b_36_57126;
  wire seg_15_4_sp4_v_b_44_57134;
  wire seg_15_4_sp4_v_b_4_56757;
  wire seg_15_4_sp4_v_t_37_57250;
  wire seg_15_5_glb_netwk_0_5;
  wire seg_15_5_glb_netwk_4_9;
  wire seg_15_5_local_g0_0_60973;
  wire seg_15_5_local_g0_5_60978;
  wire seg_15_5_local_g1_1_60982;
  wire seg_15_5_local_g1_2_60983;
  wire seg_15_5_local_g1_7_60988;
  wire seg_15_5_local_g2_2_60991;
  wire seg_15_5_local_g2_4_60993;
  wire seg_15_5_local_g3_1_60998;
  wire seg_15_5_local_g3_4_61001;
  wire seg_15_5_neigh_op_bnl_2_53151;
  wire seg_15_5_sp12_v_b_4_60411;
  wire seg_15_5_sp4_h_l_39_45749;
  wire seg_15_5_sp4_h_l_41_45751;
  wire seg_15_5_sp4_h_l_47_45747;
  wire seg_15_5_sp4_h_r_16_57244;
  wire seg_15_5_sp4_h_r_1_61068;
  wire seg_15_5_sp4_h_r_24_53407;
  wire seg_15_5_sp4_h_r_26_53411;
  wire seg_15_5_sp4_h_r_28_53413;
  wire seg_15_5_sp4_h_r_2_61071;
  wire seg_15_5_sp4_h_r_30_53415;
  wire seg_15_5_sp4_h_r_36_49577;
  wire seg_15_5_sp4_h_r_41_49582;
  wire seg_15_5_sp4_h_r_7_61076;
  wire seg_15_5_sp4_r_v_b_13_60834;
  wire seg_15_5_sp4_r_v_b_21_60842;
  wire seg_15_5_sp4_r_v_b_23_60844;
  wire seg_15_5_sp4_r_v_b_29_60960;
  wire seg_15_5_sp4_r_v_b_33_60964;
  wire seg_15_5_sp4_v_b_16_57007;
  wire seg_15_5_sp4_v_b_18_57009;
  wire seg_15_5_sp4_v_b_21_57012;
  wire seg_15_5_sp4_v_b_34_57137;
  wire seg_15_5_sp4_v_b_8_56889;
  wire seg_15_6_glb_netwk_0_5;
  wire seg_15_6_glb_netwk_4_9;
  wire seg_15_6_local_g0_0_61096;
  wire seg_15_6_local_g0_1_61097;
  wire seg_15_6_local_g0_2_61098;
  wire seg_15_6_local_g0_3_61099;
  wire seg_15_6_local_g0_4_61100;
  wire seg_15_6_local_g0_6_61102;
  wire seg_15_6_local_g1_0_61104;
  wire seg_15_6_local_g1_2_61106;
  wire seg_15_6_local_g1_3_61107;
  wire seg_15_6_local_g1_4_61108;
  wire seg_15_6_local_g1_5_61109;
  wire seg_15_6_local_g1_7_61111;
  wire seg_15_6_local_g2_0_61112;
  wire seg_15_6_local_g2_2_61114;
  wire seg_15_6_local_g2_3_61115;
  wire seg_15_6_local_g2_4_61116;
  wire seg_15_6_local_g2_5_61117;
  wire seg_15_6_local_g2_6_61118;
  wire seg_15_6_local_g3_1_61121;
  wire seg_15_6_local_g3_2_61122;
  wire seg_15_6_local_g3_3_61123;
  wire seg_15_6_local_g3_4_61124;
  wire seg_15_6_local_g3_5_61125;
  wire seg_15_6_local_g3_7_61127;
  wire seg_15_6_lutff_0_out_57225;
  wire seg_15_6_lutff_4_out_57229;
  wire seg_15_6_lutff_7_out_57232;
  wire seg_15_6_neigh_op_bnl_4_53276;
  wire seg_15_6_neigh_op_bnl_5_53277;
  wire seg_15_6_neigh_op_lft_3_53398;
  wire seg_15_6_neigh_op_lft_7_53402;
  wire seg_15_6_sp4_h_l_39_45872;
  wire seg_15_6_sp4_h_l_40_45875;
  wire seg_15_6_sp4_h_l_42_45877;
  wire seg_15_6_sp4_h_l_43_45876;
  wire seg_15_6_sp4_h_l_45_45878;
  wire seg_15_6_sp4_h_r_10_61192;
  wire seg_15_6_sp4_h_r_12_57361;
  wire seg_15_6_sp4_h_r_16_57367;
  wire seg_15_6_sp4_h_r_20_57371;
  wire seg_15_6_sp4_h_r_26_53534;
  wire seg_15_6_sp4_h_r_27_53535;
  wire seg_15_6_sp4_h_r_2_61194;
  wire seg_15_6_sp4_h_r_30_53538;
  wire seg_15_6_sp4_h_r_32_53540;
  wire seg_15_6_sp4_h_r_38_49704;
  wire seg_15_6_sp4_h_r_41_49705;
  wire seg_15_6_sp4_h_r_42_49708;
  wire seg_15_6_sp4_h_r_43_49707;
  wire seg_15_6_sp4_h_r_44_49710;
  wire seg_15_6_sp4_h_r_45_49709;
  wire seg_15_6_sp4_h_r_8_61200;
  wire seg_15_6_sp4_h_r_9_61201;
  wire seg_15_6_sp4_r_v_b_18_60962;
  wire seg_15_6_sp4_v_b_11_57013;
  wire seg_15_6_sp4_v_b_12_57126;
  wire seg_15_6_sp4_v_b_13_57127;
  wire seg_15_6_sp4_v_b_14_57128;
  wire seg_15_6_sp4_v_b_17_57131;
  wire seg_15_6_sp4_v_b_2_57006;
  wire seg_15_6_sp4_v_b_31_57255;
  wire seg_15_6_sp4_v_b_4_57008;
  wire seg_15_6_sp4_v_b_5_57007;
  wire seg_15_6_sp4_v_b_7_57009;
  wire seg_15_6_sp4_v_t_42_57501;
  wire seg_15_7_glb_netwk_0_5;
  wire seg_15_7_glb_netwk_4_9;
  wire seg_15_7_local_g1_7_61234;
  wire seg_15_7_local_g2_6_61241;
  wire seg_15_7_local_g2_7_61242;
  wire seg_15_7_local_g3_3_61246;
  wire seg_15_7_lutff_2_out_57350;
  wire seg_15_7_lutff_3_out_57351;
  wire seg_15_7_lutff_4_out_57352;
  wire seg_15_7_lutff_6_out_57354;
  wire seg_15_7_neigh_op_bot_7_57232;
  wire seg_15_7_sp12_v_b_0_60411;
  wire seg_15_7_sp4_h_l_37_45991;
  wire seg_15_7_sp4_h_l_44_46002;
  wire seg_15_7_sp4_h_l_47_45993;
  wire seg_15_7_sp4_h_r_27_53658;
  wire seg_15_7_sp4_h_r_5_61320;
  wire seg_15_7_sp4_h_r_7_61322;
  wire seg_15_7_sp4_h_r_9_61324;
  wire seg_15_7_sp4_r_v_b_15_61082;
  wire seg_15_7_sp4_v_b_10_57137;
  wire seg_15_7_sp4_v_b_9_57134;
  wire seg_15_7_sp4_v_t_36_57618;
  wire seg_15_8_glb_netwk_0_5;
  wire seg_15_8_glb_netwk_4_9;
  wire seg_15_8_local_g0_3_61345;
  wire seg_15_8_local_g0_5_61347;
  wire seg_15_8_local_g1_5_61355;
  wire seg_15_8_local_g3_0_61366;
  wire seg_15_8_lutff_2_out_57473;
  wire seg_15_8_lutff_3_out_57474;
  wire seg_15_8_lutff_4_out_57475;
  wire seg_15_8_neigh_op_lft_5_53646;
  wire seg_15_8_neigh_op_rgt_0_61301;
  wire seg_15_8_sp4_h_l_45_46124;
  wire seg_15_8_sp4_h_r_10_61438;
  wire seg_15_8_sp4_h_r_11_61439;
  wire seg_15_8_sp4_h_r_16_57613;
  wire seg_15_8_sp4_h_r_22_57609;
  wire seg_15_8_sp4_h_r_24_53776;
  wire seg_15_8_sp4_h_r_34_53778;
  wire seg_15_8_sp4_h_r_40_49952;
  wire seg_15_8_sp4_h_r_5_61443;
  wire seg_15_8_sp4_r_v_b_23_61213;
  wire seg_15_8_sp4_r_v_b_35_61335;
  wire seg_15_8_sp4_r_v_b_3_61081;
  wire seg_15_8_sp4_v_b_0_57250;
  wire seg_15_8_sp4_v_b_32_57504;
  wire seg_15_8_sp4_v_b_36_57618;
  wire seg_15_9_glb_netwk_0_5;
  wire seg_15_9_local_g0_3_61468;
  wire seg_15_9_local_g0_4_61469;
  wire seg_15_9_local_g1_2_61475;
  wire seg_15_9_local_g1_3_61476;
  wire seg_15_9_local_g2_4_61485;
  wire seg_15_9_local_g3_3_61492;
  wire seg_15_9_local_g3_7_61496;
  wire seg_15_9_neigh_op_bot_2_57473;
  wire seg_15_9_neigh_op_bot_3_57474;
  wire seg_15_9_neigh_op_bot_4_57475;
  wire seg_15_9_neigh_op_rgt_4_61428;
  wire seg_15_9_neigh_op_rgt_7_61431;
  wire seg_15_9_sp4_h_r_11_61562;
  wire seg_15_9_sp4_h_r_28_53905;
  wire seg_15_9_sp4_h_r_32_53909;
  wire seg_15_9_sp4_r_v_b_37_61572;
  wire seg_15_9_sp4_r_v_b_39_61574;
  wire seg_15_9_sp4_r_v_b_3_61204;
  wire seg_15_9_sp4_r_v_b_41_61576;
  wire seg_15_9_sp4_v_b_11_57382;
  wire seg_15_9_sp4_v_b_35_57628;
  wire seg_16_0_local_g1_3_64225;
  wire seg_16_0_span4_horz_r_0_64262;
  wire seg_16_0_span4_vert_43_60589;
  wire seg_16_10_glb_netwk_0_5;
  wire seg_16_10_glb_netwk_4_9;
  wire seg_16_10_local_g0_2_65421;
  wire seg_16_10_local_g0_4_65423;
  wire seg_16_10_local_g1_0_65427;
  wire seg_16_10_local_g1_1_65428;
  wire seg_16_10_local_g2_1_65436;
  wire seg_16_10_local_g2_3_65438;
  wire seg_16_10_local_g2_4_65439;
  wire seg_16_10_local_g3_1_65444;
  wire seg_16_10_local_g3_2_65445;
  wire seg_16_10_local_g3_3_65446;
  wire seg_16_10_lutff_1_out_61548;
  wire seg_16_10_neigh_op_rgt_1_65379;
  wire seg_16_10_neigh_op_tnl_3_57843;
  wire seg_16_10_sp4_h_l_36_50192;
  wire seg_16_10_sp4_h_l_45_50201;
  wire seg_16_10_sp4_h_l_47_50193;
  wire seg_16_10_sp4_h_r_10_65515;
  wire seg_16_10_sp4_h_r_11_65516;
  wire seg_16_10_sp4_h_r_26_57856;
  wire seg_16_10_sp4_h_r_36_54023;
  wire seg_16_10_sp4_h_r_4_65519;
  wire seg_16_10_sp4_h_r_9_65524;
  wire seg_16_10_sp4_r_v_b_17_65284;
  wire seg_16_10_sp4_r_v_b_21_65288;
  wire seg_16_10_sp4_r_v_b_23_65290;
  wire seg_16_10_sp4_r_v_b_24_65403;
  wire seg_16_10_sp4_r_v_b_29_65406;
  wire seg_16_10_sp4_r_v_b_31_65408;
  wire seg_16_10_sp4_r_v_b_33_65410;
  wire seg_16_10_sp4_r_v_b_39_65528;
  wire seg_16_10_sp4_r_v_b_41_65530;
  wire seg_16_10_sp4_r_v_b_43_65532;
  wire seg_16_10_sp4_v_b_10_61336;
  wire seg_16_10_sp4_v_b_11_61335;
  wire seg_16_10_sp4_v_b_33_61579;
  wire seg_16_10_sp4_v_b_35_61581;
  wire seg_16_10_sp4_v_b_3_61327;
  wire seg_16_10_sp4_v_b_9_61333;
  wire seg_16_10_sp4_v_t_42_61823;
  wire seg_16_11_glb_netwk_0_5;
  wire seg_16_11_glb_netwk_4_9;
  wire seg_16_11_local_g0_1_65543;
  wire seg_16_11_local_g0_2_65544;
  wire seg_16_11_local_g0_4_65546;
  wire seg_16_11_local_g0_5_65547;
  wire seg_16_11_local_g1_5_65555;
  wire seg_16_11_local_g2_4_65562;
  wire seg_16_11_local_g2_7_65565;
  wire seg_16_11_local_g3_1_65567;
  wire seg_16_11_local_g3_2_65568;
  wire seg_16_11_local_g3_3_65569;
  wire seg_16_11_local_g3_5_65571;
  wire seg_16_11_local_g3_6_65572;
  wire seg_16_11_local_g3_7_65573;
  wire seg_16_11_lutff_1_out_61671;
  wire seg_16_11_lutff_3_out_61673;
  wire seg_16_11_lutff_5_out_61675;
  wire seg_16_11_lutff_6_out_61676;
  wire seg_16_11_lutff_7_out_61677;
  wire seg_16_11_neigh_op_bnr_5_65383;
  wire seg_16_11_neigh_op_bot_1_61548;
  wire seg_16_11_neigh_op_rgt_1_65502;
  wire seg_16_11_neigh_op_rgt_2_65503;
  wire seg_16_11_neigh_op_rgt_3_65504;
  wire seg_16_11_neigh_op_rgt_4_65505;
  wire seg_16_11_neigh_op_tnl_6_57969;
  wire seg_16_11_sp12_v_b_18_65265;
  wire seg_16_11_sp12_v_b_22_65511;
  wire seg_16_11_sp4_h_l_36_50315;
  wire seg_16_11_sp4_h_l_37_50314;
  wire seg_16_11_sp4_h_l_40_50321;
  wire seg_16_11_sp4_h_l_41_50320;
  wire seg_16_11_sp4_h_r_0_65636;
  wire seg_16_11_sp4_h_r_20_61816;
  wire seg_16_11_sp4_h_r_24_57975;
  wire seg_16_11_sp4_h_r_36_54146;
  wire seg_16_11_sp4_h_r_8_65646;
  wire seg_16_11_sp4_r_v_b_21_65411;
  wire seg_16_11_sp4_r_v_b_23_65413;
  wire seg_16_11_sp4_v_b_0_61449;
  wire seg_16_11_sp4_v_b_10_61459;
  wire seg_16_11_sp4_v_b_12_61571;
  wire seg_16_11_sp4_v_b_14_61573;
  wire seg_16_11_sp4_v_b_29_61698;
  wire seg_16_11_sp4_v_b_2_61451;
  wire seg_16_11_sp4_v_b_39_61820;
  wire seg_16_11_sp4_v_b_4_61453;
  wire seg_16_12_glb_netwk_0_5;
  wire seg_16_12_local_g0_2_65667;
  wire seg_16_12_local_g0_3_65668;
  wire seg_16_12_local_g0_5_65670;
  wire seg_16_12_local_g0_7_65672;
  wire seg_16_12_local_g1_0_65673;
  wire seg_16_12_local_g1_1_65674;
  wire seg_16_12_local_g1_4_65677;
  wire seg_16_12_local_g1_5_65678;
  wire seg_16_12_local_g1_6_65679;
  wire seg_16_12_local_g1_7_65680;
  wire seg_16_12_local_g2_1_65682;
  wire seg_16_12_local_g2_5_65686;
  wire seg_16_12_local_g3_1_65690;
  wire seg_16_12_local_g3_5_65694;
  wire seg_16_12_sp4_h_l_38_50442;
  wire seg_16_12_sp4_h_l_43_50445;
  wire seg_16_12_sp4_h_l_46_50440;
  wire seg_16_12_sp4_h_r_10_65761;
  wire seg_16_12_sp4_h_r_12_61929;
  wire seg_16_12_sp4_h_r_15_61932;
  wire seg_16_12_sp4_h_r_17_61934;
  wire seg_16_12_sp4_h_r_20_61939;
  wire seg_16_12_sp4_h_r_21_61938;
  wire seg_16_12_sp4_h_r_23_61930;
  wire seg_16_12_sp4_h_r_25_58099;
  wire seg_16_12_sp4_h_r_30_58106;
  wire seg_16_12_sp4_h_r_6_65767;
  wire seg_16_12_sp4_r_v_b_45_65780;
  wire seg_16_12_sp4_v_b_0_61572;
  wire seg_16_12_sp4_v_b_13_61695;
  wire seg_16_12_sp4_v_b_19_61701;
  wire seg_16_12_sp4_v_b_37_61941;
  wire seg_16_12_sp4_v_b_41_61945;
  wire seg_16_12_sp4_v_b_4_61576;
  wire seg_16_12_sp4_v_b_5_61575;
  wire seg_16_12_sp4_v_b_6_61578;
  wire seg_16_12_sp4_v_b_7_61577;
  wire seg_16_12_sp4_v_t_40_62067;
  wire seg_16_13_glb_netwk_0_5;
  wire seg_16_13_glb_netwk_4_9;
  wire seg_16_13_local_g0_2_65790;
  wire seg_16_13_local_g0_4_65792;
  wire seg_16_13_local_g1_0_65796;
  wire seg_16_13_local_g1_1_65797;
  wire seg_16_13_local_g1_3_65799;
  wire seg_16_13_local_g1_4_65800;
  wire seg_16_13_local_g2_2_65806;
  wire seg_16_13_local_g2_3_65807;
  wire seg_16_13_local_g2_6_65810;
  wire seg_16_13_local_g3_0_65812;
  wire seg_16_13_local_g3_1_65813;
  wire seg_16_13_local_g3_2_65814;
  wire seg_16_13_local_g3_3_65815;
  wire seg_16_13_local_g3_4_65816;
  wire seg_16_13_local_g3_7_65819;
  wire seg_16_13_lutff_1_out_61917;
  wire seg_16_13_lutff_2_out_61918;
  wire seg_16_13_lutff_3_out_61919;
  wire seg_16_13_lutff_4_out_61920;
  wire seg_16_13_lutff_5_out_61921;
  wire seg_16_13_lutff_6_out_61922;
  wire seg_16_13_neigh_op_bnl_2_57965;
  wire seg_16_13_neigh_op_bnl_3_57966;
  wire seg_16_13_neigh_op_bnl_4_57967;
  wire seg_16_13_sp12_v_b_11_65020;
  wire seg_16_13_sp4_h_l_40_50567;
  wire seg_16_13_sp4_h_r_10_65884;
  wire seg_16_13_sp4_h_r_12_62052;
  wire seg_16_13_sp4_h_r_16_62058;
  wire seg_16_13_sp4_h_r_20_62062;
  wire seg_16_13_sp4_h_r_24_58221;
  wire seg_16_13_sp4_h_r_34_58223;
  wire seg_16_13_sp4_h_r_3_65887;
  wire seg_16_13_sp4_r_v_b_15_65651;
  wire seg_16_13_sp4_r_v_b_31_65777;
  wire seg_16_13_sp4_v_b_2_61697;
  wire seg_16_13_sp4_v_b_33_61948;
  wire seg_16_13_sp4_v_b_39_62066;
  wire seg_16_13_sp4_v_b_46_62073;
  wire seg_16_13_sp4_v_b_9_61702;
  wire seg_16_13_sp4_v_t_43_62193;
  wire seg_16_13_sp4_v_t_44_62194;
  wire seg_16_13_sp4_v_t_47_62197;
  wire seg_16_14_local_g0_0_65911;
  wire seg_16_14_local_g0_1_65912;
  wire seg_16_14_local_g0_2_65913;
  wire seg_16_14_local_g0_6_65917;
  wire seg_16_14_local_g1_0_65919;
  wire seg_16_14_local_g1_4_65923;
  wire seg_16_14_local_g1_5_65924;
  wire seg_16_14_local_g1_6_65925;
  wire seg_16_14_local_g1_7_65926;
  wire seg_16_14_local_g2_3_65930;
  wire seg_16_14_local_g2_6_65933;
  wire seg_16_14_local_g2_7_65934;
  wire seg_16_14_local_g3_0_65935;
  wire seg_16_14_local_g3_2_65937;
  wire seg_16_14_local_g3_3_65938;
  wire seg_16_14_local_g3_5_65940;
  wire seg_16_14_lutff_1_out_62040;
  wire seg_16_14_lutff_2_out_62041;
  wire seg_16_14_lutff_3_out_62042;
  wire seg_16_14_lutff_4_out_62043;
  wire seg_16_14_lutff_5_out_62044;
  wire seg_16_14_lutff_6_out_62045;
  wire seg_16_14_lutff_7_out_62046;
  wire seg_16_14_neigh_op_rgt_5_65875;
  wire seg_16_14_neigh_op_tnl_3_58335;
  wire seg_16_14_neigh_op_tnr_0_65993;
  wire seg_16_14_neigh_op_tnr_2_65995;
  wire seg_16_14_neigh_op_tnr_3_65996;
  wire seg_16_14_neigh_op_tnr_7_66000;
  wire seg_16_14_neigh_op_top_1_62163;
  wire seg_16_14_neigh_op_top_2_62164;
  wire seg_16_14_neigh_op_top_7_62169;
  wire seg_16_14_sp4_h_l_42_50692;
  wire seg_16_14_sp4_h_l_43_50691;
  wire seg_16_14_sp4_h_l_46_50686;
  wire seg_16_14_sp4_h_r_12_62175;
  wire seg_16_14_sp4_h_r_13_62174;
  wire seg_16_14_sp4_h_r_14_62179;
  wire seg_16_14_sp4_h_r_16_62181;
  wire seg_16_14_sp4_h_r_30_58352;
  wire seg_16_14_sp4_h_r_6_66013;
  wire seg_16_14_sp4_h_r_8_66015;
  wire seg_16_14_sp4_v_b_0_61818;
  wire seg_16_14_sp4_v_b_8_61826;
  wire seg_16_15_glb_netwk_0_5;
  wire seg_16_15_glb_netwk_4_9;
  wire seg_16_15_local_g0_6_66040;
  wire seg_16_15_local_g0_7_66041;
  wire seg_16_15_local_g1_7_66049;
  wire seg_16_15_local_g2_0_66050;
  wire seg_16_15_local_g2_1_66051;
  wire seg_16_15_local_g2_4_66054;
  wire seg_16_15_local_g3_5_66063;
  wire seg_16_15_local_g3_6_66064;
  wire seg_16_15_lutff_0_out_62162;
  wire seg_16_15_lutff_1_out_62163;
  wire seg_16_15_lutff_2_out_62164;
  wire seg_16_15_lutff_4_out_62166;
  wire seg_16_15_lutff_5_out_62167;
  wire seg_16_15_lutff_6_out_62168;
  wire seg_16_15_lutff_7_out_62169;
  wire seg_16_15_neigh_op_bnr_7_65877;
  wire seg_16_15_neigh_op_rgt_1_65994;
  wire seg_16_15_neigh_op_rgt_5_65998;
  wire seg_16_15_neigh_op_rgt_6_65999;
  wire seg_16_15_neigh_op_top_7_62292;
  wire seg_16_15_sp4_h_l_37_50806;
  wire seg_16_15_sp4_h_l_41_50812;
  wire seg_16_15_sp4_h_r_10_66130;
  wire seg_16_15_sp4_h_r_12_62298;
  wire seg_16_15_sp4_h_r_24_58467;
  wire seg_16_15_sp4_r_v_b_11_65781;
  wire seg_16_15_sp4_v_b_14_62065;
  wire seg_16_15_sp4_v_b_1_61940;
  wire seg_16_15_sp4_v_b_22_62073;
  wire seg_16_15_sp4_v_b_24_62187;
  wire seg_16_15_sp4_v_b_5_61944;
  wire seg_16_15_sp4_v_b_7_61946;
  wire seg_16_16_glb_netwk_0_5;
  wire seg_16_16_glb_netwk_1_6;
  wire seg_16_16_glb_netwk_4_9;
  wire seg_16_16_local_g0_3_66160;
  wire seg_16_16_local_g0_4_66161;
  wire seg_16_16_local_g0_5_66162;
  wire seg_16_16_local_g0_7_66164;
  wire seg_16_16_local_g1_0_66165;
  wire seg_16_16_local_g1_2_66167;
  wire seg_16_16_local_g1_4_66169;
  wire seg_16_16_local_g1_6_66171;
  wire seg_16_16_local_g1_7_66172;
  wire seg_16_16_local_g2_3_66176;
  wire seg_16_16_local_g2_7_66180;
  wire seg_16_16_local_g3_4_66185;
  wire seg_16_16_local_g3_6_66187;
  wire seg_16_16_local_g3_7_66188;
  wire seg_16_16_lutff_0_out_62285;
  wire seg_16_16_lutff_1_out_62286;
  wire seg_16_16_lutff_2_out_62287;
  wire seg_16_16_lutff_3_out_62288;
  wire seg_16_16_lutff_4_out_62289;
  wire seg_16_16_lutff_6_out_62291;
  wire seg_16_16_lutff_7_out_62292;
  wire seg_16_16_neigh_op_lft_2_58457;
  wire seg_16_16_neigh_op_lft_4_58459;
  wire seg_16_16_neigh_op_lft_5_58460;
  wire seg_16_16_neigh_op_lft_7_58462;
  wire seg_16_16_neigh_op_top_0_62408;
  wire seg_16_16_sp4_h_l_37_50929;
  wire seg_16_16_sp4_h_l_46_50932;
  wire seg_16_16_sp4_h_r_10_66253;
  wire seg_16_16_sp4_h_r_22_62423;
  wire seg_16_16_sp4_h_r_28_58596;
  wire seg_16_16_sp4_h_r_32_58600;
  wire seg_16_16_sp4_h_r_34_58592;
  wire seg_16_16_sp4_h_r_38_54765;
  wire seg_16_16_sp4_h_r_3_66256;
  wire seg_16_16_sp4_h_r_44_54771;
  wire seg_16_16_sp4_h_r_8_66261;
  wire seg_16_16_sp4_r_v_b_11_65904;
  wire seg_16_16_sp4_r_v_b_7_65900;
  wire seg_16_16_sp4_v_b_31_62315;
  wire seg_16_16_sp4_v_b_4_62068;
  wire seg_16_16_sp4_v_t_36_62555;
  wire seg_16_17_glb_netwk_0_5;
  wire seg_16_17_glb_netwk_1_6;
  wire seg_16_17_glb_netwk_4_9;
  wire seg_16_17_local_g0_0_66280;
  wire seg_16_17_local_g0_2_66282;
  wire seg_16_17_local_g0_3_66283;
  wire seg_16_17_local_g0_4_66284;
  wire seg_16_17_local_g1_5_66293;
  wire seg_16_17_local_g2_1_66297;
  wire seg_16_17_local_g2_3_66299;
  wire seg_16_17_local_g2_6_66302;
  wire seg_16_17_local_g2_7_66303;
  wire seg_16_17_local_g3_0_66304;
  wire seg_16_17_local_g3_1_66305;
  wire seg_16_17_local_g3_4_66308;
  wire seg_16_17_local_g3_6_66310;
  wire seg_16_17_lutff_0_out_62408;
  wire seg_16_17_lutff_1_out_62409;
  wire seg_16_17_lutff_2_out_62410;
  wire seg_16_17_lutff_3_out_62411;
  wire seg_16_17_lutff_4_out_62412;
  wire seg_16_17_lutff_5_out_62413;
  wire seg_16_17_lutff_6_out_62414;
  wire seg_16_17_neigh_op_bnl_1_58456;
  wire seg_16_17_neigh_op_lft_0_58578;
  wire seg_16_17_neigh_op_lft_4_58582;
  wire seg_16_17_neigh_op_tnr_6_66368;
  wire seg_16_17_sp12_v_b_0_64897;
  wire seg_16_17_sp4_h_l_38_51057;
  wire seg_16_17_sp4_h_r_14_62548;
  wire seg_16_17_sp4_h_r_19_62551;
  wire seg_16_17_sp4_h_r_24_58713;
  wire seg_16_17_sp4_h_r_38_54888;
  wire seg_16_17_sp4_h_r_3_66379;
  wire seg_16_17_sp4_r_v_b_13_66141;
  wire seg_16_17_sp4_r_v_b_15_66143;
  wire seg_16_17_sp4_r_v_b_3_66019;
  wire seg_16_17_sp4_r_v_b_43_66393;
  wire seg_16_17_sp4_r_v_b_9_66025;
  wire seg_16_17_sp4_v_b_0_62187;
  wire seg_16_17_sp4_v_b_18_62315;
  wire seg_16_17_sp4_v_b_36_62555;
  wire seg_16_17_sp4_v_b_6_62193;
  wire seg_16_18_glb_netwk_0_5;
  wire seg_16_18_glb_netwk_4_9;
  wire seg_16_18_local_g1_3_66414;
  wire seg_16_18_local_g2_6_66425;
  wire seg_16_18_sp12_v_b_0_65020;
  wire seg_16_18_sp4_r_v_b_14_66265;
  wire seg_16_18_sp4_v_b_11_62319;
  wire seg_16_1_sp4_h_l_46_49051;
  wire seg_16_20_sp12_v_b_1_65265;
  wire seg_16_22_sp12_v_b_1_65511;
  wire seg_16_2_glb_netwk_0_5;
  wire seg_16_2_glb_netwk_5_10;
  wire seg_16_2_local_g0_5_64440;
  wire seg_16_2_sp4_h_l_39_49211;
  wire seg_16_2_sp4_h_r_0_64529;
  wire seg_16_2_sp4_h_r_22_60701;
  wire seg_16_2_sp4_h_r_5_64536;
  wire seg_16_2_sp4_v_t_42_60839;
  wire seg_16_2_sp4_v_t_46_60843;
  wire seg_16_2_sp4_v_t_47_60844;
  wire seg_16_31_local_g0_6_68021;
  wire seg_16_31_local_g1_2_68025;
  wire seg_16_31_span12_vert_2_66741;
  wire seg_16_31_span12_vert_6_66987;
  wire seg_16_3_glb_netwk_0_5;
  wire seg_16_3_glb_netwk_4_9;
  wire seg_16_3_local_g0_2_64560;
  wire seg_16_3_local_g0_6_64564;
  wire seg_16_3_local_g1_2_64568;
  wire seg_16_3_local_g1_3_64569;
  wire seg_16_3_local_g2_6_64580;
  wire seg_16_3_local_g3_3_64585;
  wire seg_16_3_local_g3_4_64586;
  wire seg_16_3_lutff_2_out_60688;
  wire seg_16_3_sp12_v_b_4_64260;
  wire seg_16_3_sp4_h_l_38_49335;
  wire seg_16_3_sp4_h_l_43_49338;
  wire seg_16_3_sp4_h_r_11_64655;
  wire seg_16_3_sp4_h_r_2_64656;
  wire seg_16_3_sp4_h_r_36_53162;
  wire seg_16_3_sp4_h_r_38_53166;
  wire seg_16_3_sp4_h_r_4_64658;
  wire seg_16_3_sp4_h_r_6_64660;
  wire seg_16_3_sp4_r_v_b_23_64424;
  wire seg_16_3_sp4_r_v_b_37_64665;
  wire seg_16_3_sp4_v_b_20_60590;
  wire seg_16_3_sp4_v_b_22_60592;
  wire seg_16_3_sp4_v_b_28_60715;
  wire seg_16_3_sp4_v_b_36_60833;
  wire seg_16_3_sp4_v_b_38_60835;
  wire seg_16_3_sp4_v_b_43_60840;
  wire seg_16_4_local_g0_4_64685;
  wire seg_16_4_local_g0_7_64688;
  wire seg_16_4_local_g1_3_64692;
  wire seg_16_4_local_g1_4_64693;
  wire seg_16_4_local_g1_6_64695;
  wire seg_16_4_local_g1_7_64696;
  wire seg_16_4_local_g2_0_64697;
  wire seg_16_4_local_g2_1_64698;
  wire seg_16_4_local_g2_2_64699;
  wire seg_16_4_local_g2_3_64700;
  wire seg_16_4_local_g2_4_64701;
  wire seg_16_4_local_g2_5_64702;
  wire seg_16_4_local_g2_6_64703;
  wire seg_16_4_local_g3_0_64705;
  wire seg_16_4_local_g3_6_64711;
  wire seg_16_4_local_g3_7_64712;
  wire seg_16_4_neigh_op_bnl_2_56858;
  wire seg_16_4_neigh_op_bnr_3_64520;
  wire seg_16_4_neigh_op_bnr_4_64521;
  wire seg_16_4_neigh_op_lft_7_56986;
  wire seg_16_4_neigh_op_rgt_0_64640;
  wire seg_16_4_neigh_op_rgt_1_64641;
  wire seg_16_4_neigh_op_rgt_3_64643;
  wire seg_16_4_neigh_op_rgt_4_64644;
  wire seg_16_4_neigh_op_rgt_5_64645;
  wire seg_16_4_neigh_op_rgt_6_64646;
  wire seg_16_4_neigh_op_rgt_7_64647;
  wire seg_16_4_neigh_op_tnr_0_64763;
  wire seg_16_4_neigh_op_tnr_6_64769;
  wire seg_16_4_neigh_op_top_4_60936;
  wire seg_16_4_neigh_op_top_6_60938;
  wire seg_16_4_neigh_op_top_7_60939;
  wire seg_16_4_sp4_r_v_b_27_64666;
  wire seg_16_4_sp4_r_v_b_35_64674;
  wire seg_16_4_sp4_r_v_b_41_64792;
  wire seg_16_4_sp4_r_v_b_45_64796;
  wire seg_16_4_sp4_v_b_36_60956;
  wire seg_16_4_sp4_v_b_38_60958;
  wire seg_16_4_sp4_v_b_46_60966;
  wire seg_16_4_sp4_v_b_9_60590;
  wire seg_16_4_sp4_v_t_38_61081;
  wire seg_16_4_sp4_v_t_41_61084;
  wire seg_16_4_sp4_v_t_43_61086;
  wire seg_16_5_glb_netwk_0_5;
  wire seg_16_5_glb_netwk_4_9;
  wire seg_16_5_local_g0_1_64805;
  wire seg_16_5_local_g1_0_64812;
  wire seg_16_5_local_g1_5_64817;
  wire seg_16_5_local_g2_0_64820;
  wire seg_16_5_local_g2_2_64822;
  wire seg_16_5_local_g2_3_64823;
  wire seg_16_5_local_g2_6_64826;
  wire seg_16_5_local_g3_1_64829;
  wire seg_16_5_local_g3_2_64830;
  wire seg_16_5_local_g3_6_64834;
  wire seg_16_5_local_g3_7_64835;
  wire seg_16_5_lutff_4_out_60936;
  wire seg_16_5_lutff_5_out_60937;
  wire seg_16_5_lutff_6_out_60938;
  wire seg_16_5_lutff_7_out_60939;
  wire seg_16_5_neigh_op_rgt_0_64763;
  wire seg_16_5_neigh_op_rgt_1_64764;
  wire seg_16_5_neigh_op_rgt_2_64765;
  wire seg_16_5_neigh_op_rgt_3_64766;
  wire seg_16_5_neigh_op_rgt_6_64769;
  wire seg_16_5_neigh_op_rgt_7_64770;
  wire seg_16_5_neigh_op_tnr_2_64888;
  wire seg_16_5_neigh_op_tnr_6_64892;
  wire seg_16_5_sp12_v_b_0_64260;
  wire seg_16_5_sp4_h_l_37_49576;
  wire seg_16_5_sp4_h_l_47_49578;
  wire seg_16_5_sp4_h_r_16_61074;
  wire seg_16_5_sp4_r_v_b_39_64913;
  wire seg_16_5_sp4_r_v_b_5_64545;
  wire seg_16_5_sp4_v_b_17_60838;
  wire seg_16_5_sp4_v_b_32_60965;
  wire seg_16_5_sp4_v_b_34_60967;
  wire seg_16_5_sp4_v_b_36_61079;
  wire seg_16_5_sp4_v_b_42_61085;
  wire seg_16_6_glb_netwk_0_5;
  wire seg_16_6_glb_netwk_4_9;
  wire seg_16_6_local_g0_2_64929;
  wire seg_16_6_local_g0_4_64931;
  wire seg_16_6_local_g0_5_64932;
  wire seg_16_6_local_g0_6_64933;
  wire seg_16_6_local_g1_3_64938;
  wire seg_16_6_local_g1_6_64941;
  wire seg_16_6_local_g2_3_64946;
  wire seg_16_6_local_g3_1_64952;
  wire seg_16_6_local_g3_5_64956;
  wire seg_16_6_neigh_op_bot_5_60937;
  wire seg_16_6_sp4_h_r_10_65023;
  wire seg_16_6_sp4_h_r_20_61201;
  wire seg_16_6_sp4_h_r_24_57360;
  wire seg_16_6_sp4_h_r_28_57366;
  wire seg_16_6_sp4_h_r_3_65026;
  wire seg_16_6_sp4_r_v_b_11_64674;
  wire seg_16_6_sp4_r_v_b_17_64792;
  wire seg_16_6_sp4_r_v_b_21_64796;
  wire seg_16_6_sp4_r_v_b_23_64798;
  wire seg_16_6_sp4_r_v_b_35_64920;
  wire seg_16_6_sp4_r_v_b_3_64666;
  wire seg_16_6_sp4_v_b_0_60834;
  wire seg_16_6_sp4_v_b_10_60844;
  wire seg_16_6_sp4_v_b_12_60956;
  wire seg_16_6_sp4_v_b_14_60958;
  wire seg_16_6_sp4_v_b_1_60833;
  wire seg_16_6_sp4_v_b_22_60966;
  wire seg_16_6_sp4_v_b_3_60835;
  wire seg_16_6_sp4_v_b_42_61208;
  wire seg_16_6_sp4_v_b_46_61212;
  wire seg_16_6_sp4_v_b_5_60837;
  wire seg_16_6_sp4_v_b_8_60842;
  wire seg_16_6_sp4_v_t_36_61325;
  wire seg_16_6_sp4_v_t_42_61331;
  wire seg_16_6_sp4_v_t_46_61335;
  wire seg_16_7_glb_netwk_0_5;
  wire seg_16_7_glb_netwk_4_9;
  wire seg_16_7_local_g0_0_65050;
  wire seg_16_7_local_g0_2_65052;
  wire seg_16_7_local_g0_3_65053;
  wire seg_16_7_local_g0_4_65054;
  wire seg_16_7_local_g1_4_65062;
  wire seg_16_7_local_g1_7_65065;
  wire seg_16_7_local_g2_4_65070;
  wire seg_16_7_local_g2_7_65073;
  wire seg_16_7_lutff_3_out_61181;
  wire seg_16_7_lutff_4_out_61182;
  wire seg_16_7_neigh_op_bnr_4_64890;
  wire seg_16_7_sp4_h_l_36_49823;
  wire seg_16_7_sp4_h_l_38_49827;
  wire seg_16_7_sp4_h_r_0_65144;
  wire seg_16_7_sp4_h_r_15_61317;
  wire seg_16_7_sp4_h_r_20_61324;
  wire seg_16_7_sp4_h_r_22_61316;
  wire seg_16_7_sp4_h_r_2_65148;
  wire seg_16_7_sp4_h_r_30_57491;
  wire seg_16_7_sp4_h_r_4_65150;
  wire seg_16_7_sp4_r_v_b_13_64911;
  wire seg_16_7_sp4_r_v_b_15_64913;
  wire seg_16_7_sp4_r_v_b_29_65037;
  wire seg_16_7_sp4_r_v_b_45_65165;
  wire seg_16_7_sp4_v_b_10_60967;
  wire seg_16_7_sp4_v_b_12_61079;
  wire seg_16_7_sp4_v_b_26_61205;
  wire seg_16_7_sp4_v_b_2_60959;
  wire seg_16_7_sp4_v_b_4_60961;
  wire seg_16_7_sp4_v_b_5_60960;
  wire seg_16_7_sp4_v_b_6_60963;
  wire seg_16_7_sp4_v_b_8_60965;
  wire seg_16_7_sp4_v_b_9_60964;
  wire seg_16_7_sp4_v_t_42_61454;
  wire seg_16_8_glb_netwk_0_5;
  wire seg_16_8_glb_netwk_4_9;
  wire seg_16_8_local_g0_3_65176;
  wire seg_16_8_local_g0_7_65180;
  wire seg_16_8_local_g1_4_65185;
  wire seg_16_8_local_g1_5_65186;
  wire seg_16_8_lutff_0_out_61301;
  wire seg_16_8_sp12_h_r_3_61432;
  wire seg_16_8_sp12_h_r_5_57603;
  wire seg_16_8_sp4_h_l_37_49945;
  wire seg_16_8_sp4_h_l_45_49955;
  wire seg_16_8_sp4_h_r_20_61447;
  wire seg_16_8_sp4_h_r_2_65271;
  wire seg_16_8_sp4_h_r_4_65273;
  wire seg_16_8_sp4_h_r_8_65277;
  wire seg_16_8_sp4_v_b_34_61336;
  wire seg_16_8_sp4_v_b_40_61452;
  wire seg_16_8_sp4_v_b_5_61083;
  wire seg_16_8_sp4_v_b_7_61085;
  wire seg_16_8_sp4_v_t_36_61571;
  wire seg_16_8_sp4_v_t_38_61573;
  wire seg_16_8_sp4_v_t_39_61574;
  wire seg_16_8_sp4_v_t_43_61578;
  wire seg_16_9_glb_netwk_0_5;
  wire seg_16_9_glb_netwk_4_9;
  wire seg_16_9_local_g0_7_65303;
  wire seg_16_9_local_g1_0_65304;
  wire seg_16_9_local_g1_3_65307;
  wire seg_16_9_local_g1_6_65310;
  wire seg_16_9_local_g2_7_65319;
  wire seg_16_9_local_g3_7_65327;
  wire seg_16_9_lutff_4_out_61428;
  wire seg_16_9_lutff_7_out_61431;
  wire seg_16_9_neigh_op_rgt_7_65262;
  wire seg_16_9_sp12_h_r_12_42402;
  wire seg_16_9_sp4_h_r_11_65393;
  wire seg_16_9_sp4_h_r_24_57729;
  wire seg_16_9_sp4_h_r_34_57731;
  wire seg_16_9_sp4_h_r_42_53908;
  wire seg_16_9_sp4_h_r_46_53902;
  wire seg_16_9_sp4_r_v_b_0_65034;
  wire seg_16_9_sp4_r_v_b_15_65159;
  wire seg_16_9_sp4_r_v_b_25_65279;
  wire seg_16_9_sp4_r_v_b_6_65040;
  wire seg_16_9_sp4_v_b_10_61213;
  wire seg_16_9_sp4_v_b_11_61212;
  wire seg_16_9_sp4_v_b_12_61325;
  wire seg_16_9_sp4_v_b_2_61205;
  wire seg_16_9_sp4_v_b_34_61459;
  wire seg_16_9_sp4_v_b_3_61204;
  wire seg_16_9_sp4_v_b_42_61577;
  wire seg_16_9_sp4_v_b_7_61208;
  wire seg_17_0_span4_horz_r_12_56601;
  wire seg_17_0_span4_vert_32_64408;
  wire seg_17_10_glb_netwk_0_5;
  wire seg_17_10_glb_netwk_4_9;
  wire seg_17_10_local_g0_4_69254;
  wire seg_17_10_local_g1_0_69258;
  wire seg_17_10_local_g1_5_69263;
  wire seg_17_10_local_g1_7_69265;
  wire seg_17_10_local_g2_3_69269;
  wire seg_17_10_local_g2_4_69270;
  wire seg_17_10_local_g3_6_69280;
  wire seg_17_10_lutff_0_out_65378;
  wire seg_17_10_lutff_1_out_65379;
  wire seg_17_10_lutff_2_out_65380;
  wire seg_17_10_lutff_5_out_65383;
  wire seg_17_10_lutff_7_out_65385;
  wire seg_17_10_neigh_op_rgt_3_69212;
  wire seg_17_10_neigh_op_rgt_6_69215;
  wire seg_17_10_sp12_h_r_14_42526;
  wire seg_17_10_sp4_h_l_38_54027;
  wire seg_17_10_sp4_h_l_40_54029;
  wire seg_17_10_sp4_h_l_41_54028;
  wire seg_17_10_sp4_h_l_42_54031;
  wire seg_17_10_sp4_h_l_43_54030;
  wire seg_17_10_sp4_h_l_44_54033;
  wire seg_17_10_sp4_h_l_46_54025;
  wire seg_17_10_sp4_h_r_0_69344;
  wire seg_17_10_sp4_h_r_21_65523;
  wire seg_17_10_sp4_h_r_24_61682;
  wire seg_17_10_sp4_h_r_26_61686;
  wire seg_17_10_sp4_h_r_2_69348;
  wire seg_17_10_sp4_h_r_4_69350;
  wire seg_17_10_sp4_h_r_6_69352;
  wire seg_17_10_sp4_r_v_b_11_68997;
  wire seg_17_10_sp4_v_b_10_65167;
  wire seg_17_10_sp4_v_b_26_65405;
  wire seg_17_10_sp4_v_b_28_65407;
  wire seg_17_10_sp4_v_b_8_65165;
  wire seg_17_10_sp4_v_t_46_65658;
  wire seg_17_11_glb_netwk_0_5;
  wire seg_17_11_glb_netwk_4_9;
  wire seg_17_11_local_g0_0_69373;
  wire seg_17_11_local_g0_1_69374;
  wire seg_17_11_local_g0_5_69378;
  wire seg_17_11_local_g0_7_69380;
  wire seg_17_11_local_g1_0_69381;
  wire seg_17_11_local_g1_3_69384;
  wire seg_17_11_local_g1_4_69385;
  wire seg_17_11_local_g1_5_69386;
  wire seg_17_11_local_g1_7_69388;
  wire seg_17_11_local_g2_0_69389;
  wire seg_17_11_local_g2_2_69391;
  wire seg_17_11_local_g2_6_69395;
  wire seg_17_11_local_g3_0_69397;
  wire seg_17_11_local_g3_2_69399;
  wire seg_17_11_local_g3_5_69402;
  wire seg_17_11_local_g3_6_69403;
  wire seg_17_11_lutff_1_out_65502;
  wire seg_17_11_lutff_2_out_65503;
  wire seg_17_11_lutff_3_out_65504;
  wire seg_17_11_lutff_4_out_65505;
  wire seg_17_11_lutff_5_out_65506;
  wire seg_17_11_lutff_6_out_65507;
  wire seg_17_11_lutff_7_out_65508;
  wire seg_17_11_neigh_op_bot_0_65378;
  wire seg_17_11_neigh_op_bot_1_65379;
  wire seg_17_11_neigh_op_bot_5_65383;
  wire seg_17_11_neigh_op_lft_5_61675;
  wire seg_17_11_neigh_op_rgt_0_69332;
  wire seg_17_11_neigh_op_rgt_2_69334;
  wire seg_17_11_neigh_op_tnr_0_69455;
  wire seg_17_11_neigh_op_tnr_2_69457;
  wire seg_17_11_neigh_op_tnr_6_69461;
  wire seg_17_11_neigh_op_top_0_65624;
  wire seg_17_11_neigh_op_top_4_65628;
  wire seg_17_11_neigh_op_top_7_65631;
  wire seg_17_11_sp12_v_b_14_68850;
  wire seg_17_11_sp4_h_l_36_54146;
  wire seg_17_11_sp4_h_l_45_54155;
  wire seg_17_11_sp4_h_r_46_57978;
  wire seg_17_11_sp4_v_b_10_65290;
  wire seg_17_11_sp4_v_b_12_65402;
  wire seg_17_11_sp4_v_b_19_65409;
  wire seg_17_11_sp4_v_b_1_65279;
  wire seg_17_11_sp4_v_b_23_65413;
  wire seg_17_11_sp4_v_b_3_65281;
  wire seg_17_11_sp4_v_b_4_65284;
  wire seg_17_11_sp4_v_b_8_65288;
  wire seg_17_11_sp4_v_b_9_65287;
  wire seg_17_11_sp4_v_t_42_65777;
  wire seg_17_12_glb_netwk_0_5;
  wire seg_17_12_glb_netwk_4_9;
  wire seg_17_12_local_g0_3_69499;
  wire seg_17_12_local_g1_5_69509;
  wire seg_17_12_local_g2_3_69515;
  wire seg_17_12_local_g2_6_69518;
  wire seg_17_12_local_g3_1_69521;
  wire seg_17_12_local_g3_2_69522;
  wire seg_17_12_local_g3_5_69525;
  wire seg_17_12_local_g3_6_69526;
  wire seg_17_12_lutff_0_out_65624;
  wire seg_17_12_lutff_1_out_65625;
  wire seg_17_12_lutff_2_out_65626;
  wire seg_17_12_lutff_3_out_65627;
  wire seg_17_12_lutff_4_out_65628;
  wire seg_17_12_lutff_5_out_65629;
  wire seg_17_12_lutff_6_out_65630;
  wire seg_17_12_lutff_7_out_65631;
  wire seg_17_12_neigh_op_bnl_1_61671;
  wire seg_17_12_neigh_op_bnl_3_61673;
  wire seg_17_12_sp4_r_v_b_5_69237;
  wire seg_17_12_sp4_v_b_3_65404;
  wire seg_17_12_sp4_v_b_46_65781;
  wire seg_17_12_sp4_v_b_5_65406;
  wire seg_17_12_sp4_v_b_7_65408;
  wire seg_17_12_sp4_v_b_8_65411;
  wire seg_17_12_sp4_v_b_9_65410;
  wire seg_17_12_sp4_v_t_36_65894;
  wire seg_17_13_local_g0_4_69623;
  wire seg_17_13_local_g2_2_69637;
  wire seg_17_13_local_g2_3_69638;
  wire seg_17_13_local_g2_4_69639;
  wire seg_17_13_local_g2_6_69641;
  wire seg_17_13_local_g3_1_69644;
  wire seg_17_13_local_g3_3_69646;
  wire seg_17_13_local_g3_5_69648;
  wire seg_17_13_local_g3_7_69650;
  wire seg_17_13_lutff_2_out_65749;
  wire seg_17_13_lutff_3_out_65750;
  wire seg_17_13_lutff_4_out_65751;
  wire seg_17_13_lutff_5_out_65752;
  wire seg_17_13_lutff_6_out_65753;
  wire seg_17_13_neigh_op_tnl_1_62040;
  wire seg_17_13_neigh_op_tnl_2_62041;
  wire seg_17_13_neigh_op_tnl_3_62042;
  wire seg_17_13_neigh_op_tnl_4_62043;
  wire seg_17_13_neigh_op_tnl_5_62044;
  wire seg_17_13_neigh_op_tnl_6_62045;
  wire seg_17_13_neigh_op_tnl_7_62046;
  wire seg_17_13_neigh_op_top_4_65874;
  wire seg_17_13_sp4_h_l_39_54395;
  wire seg_17_13_sp4_h_l_45_54401;
  wire seg_17_13_sp4_h_r_27_62056;
  wire seg_17_13_sp4_h_r_2_69717;
  wire seg_17_13_sp4_v_b_2_65528;
  wire seg_17_13_sp4_v_b_4_65530;
  wire seg_17_13_sp4_v_b_6_65532;
  wire seg_17_13_sp4_v_b_8_65534;
  wire seg_17_14_glb_netwk_0_5;
  wire seg_17_14_glb_netwk_1_6;
  wire seg_17_14_glb_netwk_4_9;
  wire seg_17_14_local_g0_2_69744;
  wire seg_17_14_local_g0_4_69746;
  wire seg_17_14_local_g0_5_69747;
  wire seg_17_14_local_g0_6_69748;
  wire seg_17_14_local_g1_3_69753;
  wire seg_17_14_local_g1_4_69754;
  wire seg_17_14_local_g1_5_69755;
  wire seg_17_14_local_g1_6_69756;
  wire seg_17_14_local_g1_7_69757;
  wire seg_17_14_local_g2_0_69758;
  wire seg_17_14_local_g2_2_69760;
  wire seg_17_14_local_g2_4_69762;
  wire seg_17_14_local_g2_5_69763;
  wire seg_17_14_local_g2_6_69764;
  wire seg_17_14_local_g2_7_69765;
  wire seg_17_14_local_g3_0_69766;
  wire seg_17_14_local_g3_2_69768;
  wire seg_17_14_local_g3_4_69770;
  wire seg_17_14_local_g3_6_69772;
  wire seg_17_14_local_g3_7_69773;
  wire seg_17_14_lutff_1_out_65871;
  wire seg_17_14_lutff_2_out_65872;
  wire seg_17_14_lutff_3_out_65873;
  wire seg_17_14_lutff_4_out_65874;
  wire seg_17_14_lutff_5_out_65875;
  wire seg_17_14_lutff_6_out_65876;
  wire seg_17_14_lutff_7_out_65877;
  wire seg_17_14_neigh_op_bot_2_65749;
  wire seg_17_14_neigh_op_bot_3_65750;
  wire seg_17_14_neigh_op_bot_4_65751;
  wire seg_17_14_neigh_op_bot_5_65752;
  wire seg_17_14_neigh_op_bot_6_65753;
  wire seg_17_14_neigh_op_tnl_0_62162;
  wire seg_17_14_neigh_op_top_4_65997;
  wire seg_17_14_neigh_op_top_7_66000;
  wire seg_17_14_sp4_h_l_39_54518;
  wire seg_17_14_sp4_h_r_0_69836;
  wire seg_17_14_sp4_h_r_14_66010;
  wire seg_17_14_sp4_h_r_30_62182;
  wire seg_17_14_sp4_h_r_34_62176;
  wire seg_17_14_sp4_h_r_3_69841;
  wire seg_17_14_sp4_h_r_5_69843;
  wire seg_17_14_sp4_v_b_28_65899;
  wire seg_17_14_sp4_v_b_2_65651;
  wire seg_17_14_sp4_v_b_30_65901;
  wire seg_17_14_sp4_v_b_31_65900;
  wire seg_17_14_sp4_v_b_32_65903;
  wire seg_17_14_sp4_v_b_34_65905;
  wire seg_17_14_sp4_v_b_36_66017;
  wire seg_17_14_sp4_v_b_40_66021;
  wire seg_17_14_sp4_v_t_38_66142;
  wire seg_17_15_glb_netwk_0_5;
  wire seg_17_15_glb_netwk_4_9;
  wire seg_17_15_local_g0_3_69868;
  wire seg_17_15_local_g2_1_69882;
  wire seg_17_15_local_g2_2_69883;
  wire seg_17_15_local_g2_3_69884;
  wire seg_17_15_local_g2_5_69886;
  wire seg_17_15_local_g3_2_69891;
  wire seg_17_15_local_g3_3_69892;
  wire seg_17_15_local_g3_5_69894;
  wire seg_17_15_lutff_0_out_65993;
  wire seg_17_15_lutff_1_out_65994;
  wire seg_17_15_lutff_2_out_65995;
  wire seg_17_15_lutff_3_out_65996;
  wire seg_17_15_lutff_4_out_65997;
  wire seg_17_15_lutff_5_out_65998;
  wire seg_17_15_lutff_6_out_65999;
  wire seg_17_15_lutff_7_out_66000;
  wire seg_17_15_neigh_op_tnl_2_62287;
  wire seg_17_15_neigh_op_tnl_3_62288;
  wire seg_17_15_neigh_op_tnr_2_69949;
  wire seg_17_15_neigh_op_tnr_5_69952;
  wire seg_17_15_sp4_h_r_4_69965;
  wire seg_17_15_sp4_r_v_b_27_69850;
  wire seg_17_15_sp4_r_v_b_3_69604;
  wire seg_17_15_sp4_r_v_b_9_69610;
  wire seg_17_15_sp4_v_b_12_65894;
  wire seg_17_15_sp4_v_b_1_65771;
  wire seg_17_15_sp4_v_b_27_66019;
  wire seg_17_15_sp4_v_b_33_66025;
  wire seg_17_15_sp4_v_b_37_66141;
  wire seg_17_15_sp4_v_b_3_65773;
  wire seg_17_15_sp4_v_b_7_65777;
  wire seg_17_16_local_g0_2_69990;
  wire seg_17_16_local_g0_3_69991;
  wire seg_17_16_local_g1_1_69997;
  wire seg_17_16_local_g1_4_70000;
  wire seg_17_16_local_g1_5_70001;
  wire seg_17_16_local_g1_6_70002;
  wire seg_17_16_local_g1_7_70003;
  wire seg_17_16_local_g2_4_70008;
  wire seg_17_16_local_g3_4_70016;
  wire seg_17_16_lutff_1_out_66117;
  wire seg_17_16_neigh_op_bnr_1_69825;
  wire seg_17_16_neigh_op_bnr_2_69826;
  wire seg_17_16_neigh_op_bnr_3_69827;
  wire seg_17_16_neigh_op_bnr_4_69828;
  wire seg_17_16_neigh_op_bnr_5_69829;
  wire seg_17_16_neigh_op_bnr_6_69830;
  wire seg_17_16_neigh_op_bnr_7_69831;
  wire seg_17_16_neigh_op_rgt_4_69951;
  wire seg_17_16_neigh_op_tnr_4_70074;
  wire seg_17_16_sp4_v_b_10_65905;
  wire seg_17_16_sp4_v_b_11_65904;
  wire seg_17_16_sp4_v_b_12_66017;
  wire seg_17_16_sp4_v_b_3_65896;
  wire seg_17_16_sp4_v_b_4_65899;
  wire seg_17_16_sp4_v_b_6_65901;
  wire seg_17_16_sp4_v_b_8_65903;
  wire seg_17_16_sp4_v_t_41_66391;
  wire seg_17_16_sp4_v_t_43_66393;
  wire seg_17_17_glb_netwk_0_5;
  wire seg_17_17_glb_netwk_1_6;
  wire seg_17_17_glb_netwk_4_9;
  wire seg_17_17_local_g0_0_70111;
  wire seg_17_17_local_g0_3_70114;
  wire seg_17_17_local_g0_4_70115;
  wire seg_17_17_local_g0_5_70116;
  wire seg_17_17_local_g0_6_70117;
  wire seg_17_17_local_g0_7_70118;
  wire seg_17_17_local_g1_0_70119;
  wire seg_17_17_local_g1_1_70120;
  wire seg_17_17_local_g1_5_70124;
  wire seg_17_17_local_g2_4_70131;
  wire seg_17_17_local_g2_7_70134;
  wire seg_17_17_local_g3_3_70138;
  wire seg_17_17_lutff_0_out_66239;
  wire seg_17_17_lutff_3_out_66242;
  wire seg_17_17_lutff_4_out_66243;
  wire seg_17_17_lutff_5_out_66244;
  wire seg_17_17_neigh_op_bnr_0_69947;
  wire seg_17_17_neigh_op_bnr_4_69951;
  wire seg_17_17_neigh_op_bot_1_66117;
  wire seg_17_17_neigh_op_rgt_4_70074;
  wire seg_17_17_neigh_op_top_6_66368;
  wire seg_17_17_sp4_h_r_14_66379;
  wire seg_17_17_sp4_h_r_24_62543;
  wire seg_17_17_sp4_h_r_39_58717;
  wire seg_17_17_sp4_h_r_40_58720;
  wire seg_17_17_sp4_h_r_46_58716;
  wire seg_17_17_sp4_r_v_b_13_69972;
  wire seg_17_17_sp4_r_v_b_3_69850;
  wire seg_17_17_sp4_v_b_11_66027;
  wire seg_17_17_sp4_v_b_14_66142;
  wire seg_17_17_sp4_v_b_15_66143;
  wire seg_17_17_sp4_v_b_19_66147;
  wire seg_17_17_sp4_v_b_5_66021;
  wire seg_17_17_sp4_v_b_8_66026;
  wire seg_17_18_glb_netwk_0_5;
  wire seg_17_18_glb_netwk_4_9;
  wire seg_17_18_local_g0_4_70238;
  wire seg_17_18_lutff_6_out_66368;
  wire seg_17_18_neigh_op_bot_4_66243;
  wire seg_17_18_sp12_v_b_1_68850;
  wire seg_17_18_sp4_h_r_44_58847;
  wire seg_17_18_sp4_v_b_28_66391;
  wire seg_17_19_sp4_v_b_1_66263;
  wire seg_17_23_sp4_v_b_4_66760;
  wire seg_17_27_sp4_v_b_7_67253;
  wire seg_17_2_glb_netwk_0_5;
  wire seg_17_2_glb_netwk_5_10;
  wire seg_17_2_local_g1_7_68281;
  wire seg_17_2_local_g3_2_68292;
  wire seg_17_2_sp4_h_r_0_68360;
  wire seg_17_2_sp4_h_r_14_64534;
  wire seg_17_2_sp4_r_v_b_18_68238;
  wire seg_17_2_sp4_v_b_15_64401;
  wire seg_17_30_sp12_v_b_1_70326;
  wire seg_17_31_local_g1_1_71855;
  wire seg_17_31_span4_vert_1_67739;
  wire seg_17_31_span4_vert_7_67745;
  wire seg_17_3_glb_netwk_0_5;
  wire seg_17_3_glb_netwk_4_9;
  wire seg_17_3_local_g0_2_68391;
  wire seg_17_3_local_g0_3_68392;
  wire seg_17_3_local_g1_3_68400;
  wire seg_17_3_local_g2_4_68409;
  wire seg_17_3_local_g3_0_68413;
  wire seg_17_3_lutff_0_out_64517;
  wire seg_17_3_lutff_1_out_64518;
  wire seg_17_3_lutff_3_out_64520;
  wire seg_17_3_lutff_4_out_64521;
  wire seg_17_3_sp4_h_l_39_53165;
  wire seg_17_3_sp4_h_l_47_53163;
  wire seg_17_3_sp4_h_r_10_68485;
  wire seg_17_3_sp4_h_r_11_68486;
  wire seg_17_3_sp4_h_r_36_56992;
  wire seg_17_3_sp4_h_r_3_68488;
  wire seg_17_3_sp4_r_v_b_36_68495;
  wire seg_17_3_sp4_v_b_8_64408;
  wire seg_17_4_glb_netwk_0_5;
  wire seg_17_4_glb_netwk_4_9;
  wire seg_17_4_local_g0_3_68515;
  wire seg_17_4_local_g1_0_68520;
  wire seg_17_4_local_g1_2_68522;
  wire seg_17_4_local_g1_3_68523;
  wire seg_17_4_local_g1_5_68525;
  wire seg_17_4_local_g1_6_68526;
  wire seg_17_4_local_g1_7_68527;
  wire seg_17_4_local_g2_7_68535;
  wire seg_17_4_lutff_0_out_64640;
  wire seg_17_4_lutff_1_out_64641;
  wire seg_17_4_lutff_3_out_64643;
  wire seg_17_4_lutff_4_out_64644;
  wire seg_17_4_lutff_5_out_64645;
  wire seg_17_4_lutff_6_out_64646;
  wire seg_17_4_lutff_7_out_64647;
  wire seg_17_4_sp12_h_r_3_64771;
  wire seg_17_4_sp4_h_l_37_53284;
  wire seg_17_4_sp4_h_l_39_53288;
  wire seg_17_4_sp4_h_l_44_53295;
  wire seg_17_4_sp4_h_l_47_53286;
  wire seg_17_4_sp4_h_r_21_64785;
  wire seg_17_4_sp4_h_r_23_64777;
  wire seg_17_4_sp4_h_r_3_68611;
  wire seg_17_4_sp4_r_v_b_0_68244;
  wire seg_17_4_sp4_r_v_b_15_68375;
  wire seg_17_4_sp4_r_v_b_32_68504;
  wire seg_17_4_sp4_r_v_b_5_68248;
  wire seg_17_4_sp4_v_b_10_64424;
  wire seg_17_4_sp4_v_b_18_64547;
  wire seg_17_4_sp4_v_b_22_64551;
  wire seg_17_4_sp4_v_t_36_64910;
  wire seg_17_4_sp4_v_t_38_64912;
  wire seg_17_4_sp4_v_t_40_64914;
  wire seg_17_5_glb_netwk_0_5;
  wire seg_17_5_glb_netwk_4_9;
  wire seg_17_5_local_g0_3_68638;
  wire seg_17_5_local_g0_7_68642;
  wire seg_17_5_local_g1_0_68643;
  wire seg_17_5_local_g1_1_68644;
  wire seg_17_5_local_g1_3_68646;
  wire seg_17_5_local_g2_2_68653;
  wire seg_17_5_local_g3_7_68666;
  wire seg_17_5_lutff_0_out_64763;
  wire seg_17_5_lutff_1_out_64764;
  wire seg_17_5_lutff_2_out_64765;
  wire seg_17_5_lutff_3_out_64766;
  wire seg_17_5_lutff_5_out_64768;
  wire seg_17_5_lutff_6_out_64769;
  wire seg_17_5_lutff_7_out_64770;
  wire seg_17_5_sp4_h_l_37_53407;
  wire seg_17_5_sp4_h_l_39_53411;
  wire seg_17_5_sp4_h_l_43_53415;
  wire seg_17_5_sp4_h_r_11_68732;
  wire seg_17_5_sp4_h_r_15_64902;
  wire seg_17_5_sp4_h_r_16_64905;
  wire seg_17_5_sp4_h_r_1_68730;
  wire seg_17_5_sp4_h_r_3_68734;
  wire seg_17_5_sp4_h_r_5_68736;
  wire seg_17_5_sp4_h_r_7_68738;
  wire seg_17_5_sp4_r_v_b_10_68383;
  wire seg_17_5_sp4_r_v_b_47_68752;
  wire seg_17_5_sp4_v_t_45_65042;
  wire seg_17_6_glb_netwk_0_5;
  wire seg_17_6_glb_netwk_4_9;
  wire seg_17_6_local_g0_6_68764;
  wire seg_17_6_local_g1_5_68771;
  wire seg_17_6_local_g2_5_68779;
  wire seg_17_6_local_g3_1_68783;
  wire seg_17_6_local_g3_3_68785;
  wire seg_17_6_lutff_2_out_64888;
  wire seg_17_6_lutff_4_out_64890;
  wire seg_17_6_lutff_5_out_64891;
  wire seg_17_6_lutff_6_out_64892;
  wire seg_17_6_neigh_op_rgt_3_68720;
  wire seg_17_6_sp4_h_l_37_53530;
  wire seg_17_6_sp4_h_l_40_53537;
  wire seg_17_6_sp4_h_l_47_53532;
  wire seg_17_6_sp4_h_r_14_65026;
  wire seg_17_6_sp4_h_r_22_65024;
  wire seg_17_6_sp4_h_r_5_68859;
  wire seg_17_6_sp4_r_v_b_17_68623;
  wire seg_17_6_sp4_v_b_0_64665;
  wire seg_17_6_sp4_v_t_47_65167;
  wire seg_17_7_glb_netwk_0_5;
  wire seg_17_7_glb_netwk_4_9;
  wire seg_17_7_local_g0_7_68888;
  wire seg_17_7_local_g2_2_68899;
  wire seg_17_7_lutff_7_out_65016;
  wire seg_17_7_sp4_h_r_3_68980;
  wire seg_17_7_sp4_h_r_46_57486;
  wire seg_17_7_sp4_h_r_7_68984;
  wire seg_17_7_sp4_h_r_9_68986;
  wire seg_17_7_sp4_v_b_10_64798;
  wire seg_17_7_sp4_v_b_14_64912;
  wire seg_17_7_sp4_v_b_34_65044;
  wire seg_17_8_glb_netwk_0_5;
  wire seg_17_8_local_g0_1_69005;
  wire seg_17_8_local_g0_2_69006;
  wire seg_17_8_local_g0_5_69009;
  wire seg_17_8_local_g1_1_69013;
  wire seg_17_8_local_g1_2_69014;
  wire seg_17_8_local_g1_7_69019;
  wire seg_17_8_local_g2_0_69020;
  wire seg_17_8_local_g2_2_69022;
  wire seg_17_8_local_g2_4_69024;
  wire seg_17_8_local_g3_0_69028;
  wire seg_17_8_local_g3_2_69030;
  wire seg_17_8_local_g3_4_69032;
  wire seg_17_8_sp4_h_l_36_53777;
  wire seg_17_8_sp4_h_l_39_53780;
  wire seg_17_8_sp4_h_l_43_53784;
  wire seg_17_8_sp4_h_l_47_53778;
  wire seg_17_8_sp4_h_r_18_65276;
  wire seg_17_8_sp4_h_r_1_69099;
  wire seg_17_8_sp4_h_r_2_69102;
  wire seg_17_8_sp4_h_r_32_61446;
  wire seg_17_8_sp4_h_r_34_61438;
  wire seg_17_8_sp4_h_r_36_57607;
  wire seg_17_8_sp4_h_r_42_57615;
  wire seg_17_8_sp4_h_r_44_57617;
  wire seg_17_8_sp4_h_r_5_69105;
  wire seg_17_8_sp4_h_r_7_69107;
  wire seg_17_8_sp4_r_v_b_16_68868;
  wire seg_17_8_sp4_r_v_b_18_68870;
  wire seg_17_8_sp4_v_b_0_64911;
  wire seg_17_8_sp4_v_b_10_64921;
  wire seg_17_8_sp4_v_b_11_64920;
  wire seg_17_8_sp4_v_b_15_65036;
  wire seg_17_8_sp4_v_b_17_65038;
  wire seg_17_8_sp4_v_b_28_65161;
  wire seg_17_8_sp4_v_b_9_64918;
  wire seg_17_8_sp4_v_t_36_65402;
  wire seg_17_8_sp4_v_t_39_65405;
  wire seg_17_9_glb_netwk_0_5;
  wire seg_17_9_glb_netwk_4_9;
  wire seg_17_9_local_g0_1_69128;
  wire seg_17_9_local_g0_4_69131;
  wire seg_17_9_lutff_7_out_65262;
  wire seg_17_9_sp4_h_l_41_53905;
  wire seg_17_9_sp4_h_l_45_53909;
  wire seg_17_9_sp4_h_l_47_53901;
  wire seg_17_9_sp4_h_r_1_69222;
  wire seg_17_9_sp4_h_r_20_65401;
  wire seg_17_9_sp4_h_r_6_69229;
  wire seg_17_9_sp4_h_r_7_69230;
  wire seg_17_9_sp4_v_b_5_65037;
  wire seg_17_9_sp4_v_b_8_65042;
  wire seg_18_0_local_g1_0_71884;
  wire seg_18_0_span4_horz_r_12_60431;
  wire seg_18_0_span4_vert_24_68230;
  wire seg_18_10_glb_netwk_0_5;
  wire seg_18_10_glb_netwk_4_9;
  wire seg_18_10_local_g0_0_73081;
  wire seg_18_10_local_g0_1_73082;
  wire seg_18_10_local_g0_5_73086;
  wire seg_18_10_local_g0_6_73087;
  wire seg_18_10_local_g1_2_73091;
  wire seg_18_10_local_g1_5_73094;
  wire seg_18_10_local_g1_6_73095;
  wire seg_18_10_local_g1_7_73096;
  wire seg_18_10_local_g2_0_73097;
  wire seg_18_10_local_g2_6_73103;
  wire seg_18_10_local_g2_7_73104;
  wire seg_18_10_local_g3_1_73106;
  wire seg_18_10_local_g3_2_73107;
  wire seg_18_10_lutff_1_out_69210;
  wire seg_18_10_lutff_3_out_69212;
  wire seg_18_10_lutff_4_out_69213;
  wire seg_18_10_lutff_6_out_69215;
  wire seg_18_10_neigh_op_bot_5_69091;
  wire seg_18_10_neigh_op_bot_6_69092;
  wire seg_18_10_neigh_op_lft_2_65380;
  wire seg_18_10_neigh_op_top_7_69339;
  wire seg_18_10_sp4_h_r_0_73175;
  wire seg_18_10_sp4_h_r_16_69351;
  wire seg_18_10_sp4_h_r_21_69354;
  wire seg_18_10_sp4_h_r_26_65517;
  wire seg_18_10_sp4_h_r_30_65521;
  wire seg_18_10_sp4_h_r_40_61689;
  wire seg_18_10_sp4_h_r_42_61691;
  wire seg_18_10_sp4_h_r_5_73182;
  wire seg_18_10_sp4_r_v_b_21_72950;
  wire seg_18_10_sp4_v_b_17_69115;
  wire seg_18_10_sp4_v_b_1_68987;
  wire seg_18_10_sp4_v_b_22_69120;
  wire seg_18_10_sp4_v_b_38_69358;
  wire seg_18_10_sp4_v_b_3_68989;
  wire seg_18_10_sp4_v_b_47_69367;
  wire seg_18_10_sp4_v_b_7_68993;
  wire seg_18_10_sp4_v_b_8_68996;
  wire seg_18_10_sp4_v_b_9_68995;
  wire seg_18_11_glb_netwk_0_5;
  wire seg_18_11_glb_netwk_4_9;
  wire seg_18_11_local_g0_1_73205;
  wire seg_18_11_local_g0_6_73210;
  wire seg_18_11_local_g0_7_73211;
  wire seg_18_11_local_g1_6_73218;
  wire seg_18_11_local_g2_0_73220;
  wire seg_18_11_local_g2_3_73223;
  wire seg_18_11_local_g2_5_73225;
  wire seg_18_11_local_g3_0_73228;
  wire seg_18_11_lutff_0_out_69332;
  wire seg_18_11_lutff_1_out_69333;
  wire seg_18_11_lutff_2_out_69334;
  wire seg_18_11_lutff_3_out_69335;
  wire seg_18_11_lutff_5_out_69337;
  wire seg_18_11_lutff_6_out_69338;
  wire seg_18_11_lutff_7_out_69339;
  wire seg_18_11_neigh_op_lft_6_65507;
  wire seg_18_11_neigh_op_lft_7_65508;
  wire seg_18_11_sp4_h_l_37_57975;
  wire seg_18_11_sp4_h_r_24_65636;
  wire seg_18_11_sp4_h_r_32_65646;
  wire seg_18_11_sp4_h_r_40_61812;
  wire seg_18_11_sp4_h_r_6_73306;
  wire seg_18_11_sp4_h_r_8_73308;
  wire seg_18_11_sp4_v_b_24_69357;
  wire seg_18_11_sp4_v_b_40_69483;
  wire seg_18_11_sp4_v_t_36_69602;
  wire seg_18_12_glb_netwk_0_5;
  wire seg_18_12_glb_netwk_4_9;
  wire seg_18_12_local_g0_3_73330;
  wire seg_18_12_local_g0_4_73331;
  wire seg_18_12_local_g1_0_73335;
  wire seg_18_12_local_g1_1_73336;
  wire seg_18_12_local_g1_7_73342;
  wire seg_18_12_local_g3_1_73352;
  wire seg_18_12_local_g3_2_73353;
  wire seg_18_12_lutff_0_out_69455;
  wire seg_18_12_lutff_1_out_69456;
  wire seg_18_12_lutff_2_out_69457;
  wire seg_18_12_lutff_3_out_69458;
  wire seg_18_12_lutff_4_out_69459;
  wire seg_18_12_lutff_6_out_69461;
  wire seg_18_12_neigh_op_lft_1_65625;
  wire seg_18_12_neigh_op_top_0_69578;
  wire seg_18_12_sp4_h_r_11_73424;
  wire seg_18_12_sp4_h_r_15_69594;
  wire seg_18_12_sp4_v_b_14_69358;
  wire seg_18_12_sp4_v_b_34_69490;
  wire seg_18_12_sp4_v_b_6_69240;
  wire seg_18_12_sp4_v_t_39_69728;
  wire seg_18_13_glb_netwk_0_5;
  wire seg_18_13_glb_netwk_4_9;
  wire seg_18_13_local_g0_1_73451;
  wire seg_18_13_local_g1_1_73459;
  wire seg_18_13_local_g2_1_73467;
  wire seg_18_13_local_g3_1_73475;
  wire seg_18_13_local_g3_3_73477;
  wire seg_18_13_local_g3_7_73481;
  wire seg_18_13_lutff_0_out_69578;
  wire seg_18_13_neigh_op_top_1_69702;
  wire seg_18_13_sp4_h_r_34_65884;
  wire seg_18_13_sp4_h_r_36_62052;
  wire seg_18_13_sp4_h_r_40_62058;
  wire seg_18_13_sp4_h_r_44_62062;
  wire seg_18_13_sp4_v_b_0_69357;
  wire seg_18_13_sp4_v_b_10_69367;
  wire seg_18_13_sp4_v_b_17_69484;
  wire seg_18_13_sp4_v_b_27_69604;
  wire seg_18_13_sp4_v_b_33_69610;
  wire seg_18_13_sp4_v_b_41_69730;
  wire seg_18_13_sp4_v_b_47_69736;
  wire seg_18_13_sp4_v_b_8_69365;
  wire seg_18_14_glb_netwk_0_5;
  wire seg_18_14_glb_netwk_4_9;
  wire seg_18_14_local_g0_0_73573;
  wire seg_18_14_local_g0_2_73575;
  wire seg_18_14_local_g0_3_73576;
  wire seg_18_14_local_g1_1_73582;
  wire seg_18_14_local_g1_3_73584;
  wire seg_18_14_local_g1_6_73587;
  wire seg_18_14_local_g2_1_73590;
  wire seg_18_14_local_g3_2_73599;
  wire seg_18_14_lutff_0_out_69701;
  wire seg_18_14_lutff_1_out_69702;
  wire seg_18_14_lutff_2_out_69703;
  wire seg_18_14_lutff_3_out_69704;
  wire seg_18_14_lutff_4_out_69705;
  wire seg_18_14_lutff_7_out_69708;
  wire seg_18_14_neigh_op_lft_1_65871;
  wire seg_18_14_neigh_op_lft_2_65872;
  wire seg_18_14_neigh_op_lft_3_65873;
  wire seg_18_14_neigh_op_lft_6_65876;
  wire seg_18_14_sp4_h_l_41_58350;
  wire seg_18_14_sp4_h_l_44_58355;
  wire seg_18_14_sp4_h_l_45_58354;
  wire seg_18_14_sp4_h_l_47_58346;
  wire seg_18_14_sp4_h_r_0_73667;
  wire seg_18_14_sp4_h_r_11_73670;
  wire seg_18_14_sp4_h_r_26_66009;
  wire seg_18_14_sp4_h_r_30_66013;
  wire seg_18_14_sp4_h_r_32_66015;
  wire seg_18_14_sp4_h_r_36_62175;
  wire seg_18_14_sp4_h_r_38_62179;
  wire seg_18_14_sp4_h_r_40_62181;
  wire seg_18_14_sp4_h_r_41_62180;
  wire seg_18_14_sp4_r_v_b_11_73320;
  wire seg_18_14_sp4_v_b_12_69602;
  wire seg_18_14_sp4_v_b_3_69481;
  wire seg_18_14_sp4_v_t_37_69972;
  wire seg_18_14_sp4_v_t_43_69978;
  wire seg_18_15_local_g0_1_73697;
  wire seg_18_15_local_g0_2_73698;
  wire seg_18_15_local_g0_4_73700;
  wire seg_18_15_local_g0_5_73701;
  wire seg_18_15_local_g0_6_73702;
  wire seg_18_15_local_g0_7_73703;
  wire seg_18_15_local_g1_0_73704;
  wire seg_18_15_local_g1_1_73705;
  wire seg_18_15_local_g1_2_73706;
  wire seg_18_15_local_g1_3_73707;
  wire seg_18_15_local_g1_4_73708;
  wire seg_18_15_local_g1_5_73709;
  wire seg_18_15_local_g1_7_73711;
  wire seg_18_15_local_g3_2_73722;
  wire seg_18_15_local_g3_3_73723;
  wire seg_18_15_local_g3_4_73724;
  wire seg_18_15_lutff_1_out_69825;
  wire seg_18_15_lutff_2_out_69826;
  wire seg_18_15_lutff_3_out_69827;
  wire seg_18_15_lutff_4_out_69828;
  wire seg_18_15_lutff_5_out_69829;
  wire seg_18_15_lutff_6_out_69830;
  wire seg_18_15_lutff_7_out_69831;
  wire seg_18_15_neigh_op_bot_0_69701;
  wire seg_18_15_neigh_op_bot_2_69703;
  wire seg_18_15_neigh_op_bot_3_69704;
  wire seg_18_15_neigh_op_bot_4_69705;
  wire seg_18_15_neigh_op_bot_7_69708;
  wire seg_18_15_neigh_op_lft_1_65994;
  wire seg_18_15_neigh_op_lft_4_65997;
  wire seg_18_15_neigh_op_lft_5_65998;
  wire seg_18_15_neigh_op_lft_6_65999;
  wire seg_18_15_neigh_op_lft_7_66000;
  wire seg_18_15_neigh_op_top_2_69949;
  wire seg_18_15_neigh_op_top_5_69952;
  wire seg_18_15_sp4_h_l_37_58467;
  wire seg_18_15_sp4_h_r_17_69965;
  wire seg_18_15_sp4_h_r_34_66130;
  wire seg_18_15_sp4_h_r_36_62298;
  wire seg_18_15_sp4_v_b_43_69978;
  wire seg_18_16_glb_netwk_0_5;
  wire seg_18_16_glb_netwk_4_9;
  wire seg_18_16_local_g0_0_73819;
  wire seg_18_16_local_g1_3_73830;
  wire seg_18_16_local_g2_0_73835;
  wire seg_18_16_local_g2_4_73839;
  wire seg_18_16_local_g2_6_73841;
  wire seg_18_16_local_g3_0_73843;
  wire seg_18_16_local_g3_1_73844;
  wire seg_18_16_local_g3_5_73848;
  wire seg_18_16_local_g3_7_73850;
  wire seg_18_16_lutff_0_out_69947;
  wire seg_18_16_lutff_1_out_69948;
  wire seg_18_16_lutff_2_out_69949;
  wire seg_18_16_lutff_4_out_69951;
  wire seg_18_16_lutff_5_out_69952;
  wire seg_18_16_neigh_op_bnl_4_65997;
  wire seg_18_16_neigh_op_bnl_7_66000;
  wire seg_18_16_neigh_op_tnl_0_66239;
  wire seg_18_16_sp12_v_b_1_72435;
  wire seg_18_16_sp4_h_r_16_70089;
  wire seg_18_16_sp4_h_r_19_70090;
  wire seg_18_16_sp4_h_r_32_66261;
  wire seg_18_16_sp4_h_r_34_66253;
  wire seg_18_16_sp4_r_v_b_14_73681;
  wire seg_18_16_sp4_v_b_10_69736;
  wire seg_18_16_sp4_v_b_2_69728;
  wire seg_18_16_sp4_v_b_30_69978;
  wire seg_18_16_sp4_v_b_37_70095;
  wire seg_18_16_sp4_v_b_4_69730;
  wire seg_18_17_glb_netwk_0_5;
  wire seg_18_17_glb_netwk_4_9;
  wire seg_18_17_local_g3_7_73973;
  wire seg_18_17_lutff_4_out_70074;
  wire seg_18_17_sp4_h_r_39_62547;
  wire seg_18_18_sp4_v_b_9_69979;
  wire seg_18_22_sp4_v_b_0_70464;
  wire seg_18_26_sp4_v_b_8_70964;
  wire seg_18_2_glb_netwk_0_5;
  wire seg_18_2_glb_netwk_4_9;
  wire seg_18_2_local_g0_6_72103;
  wire seg_18_2_local_g1_4_72109;
  wire seg_18_2_local_g2_3_72116;
  wire seg_18_2_sp4_h_r_12_68361;
  wire seg_18_2_sp4_h_r_22_68363;
  wire seg_18_2_sp4_h_r_24_64529;
  wire seg_18_2_sp4_h_r_35_64532;
  wire seg_18_2_sp4_h_r_40_60705;
  wire seg_18_30_sp4_v_b_11_71457;
  wire seg_18_31_local_g0_2_75679;
  wire seg_18_31_local_g0_5_75682;
  wire seg_18_31_span4_horz_r_5_71863;
  wire seg_18_31_span4_vert_42_75661;
  wire seg_18_3_glb_netwk_0_5;
  wire seg_18_3_glb_netwk_4_9;
  wire seg_18_3_local_g0_2_72222;
  wire seg_18_3_local_g0_3_72223;
  wire seg_18_3_local_g0_4_72224;
  wire seg_18_3_local_g1_0_72228;
  wire seg_18_3_local_g1_1_72229;
  wire seg_18_3_local_g1_5_72233;
  wire seg_18_3_local_g1_7_72235;
  wire seg_18_3_local_g3_5_72249;
  wire seg_18_3_lutff_0_out_68348;
  wire seg_18_3_lutff_1_out_68349;
  wire seg_18_3_lutff_2_out_68350;
  wire seg_18_3_lutff_3_out_68351;
  wire seg_18_3_lutff_4_out_68352;
  wire seg_18_3_lutff_5_out_68353;
  wire seg_18_3_lutff_7_out_68355;
  wire seg_18_3_sp4_h_l_42_57000;
  wire seg_18_3_sp4_h_r_11_72317;
  wire seg_18_3_sp4_h_r_18_68492;
  wire seg_18_3_sp4_h_r_1_72315;
  wire seg_18_3_sp4_h_r_21_68493;
  wire seg_18_3_sp4_h_r_4_72320;
  wire seg_18_3_sp4_h_r_8_72324;
  wire seg_18_3_sp4_r_v_b_7_72069;
  wire seg_18_3_sp4_v_b_44_68503;
  wire seg_18_3_sp4_v_t_44_68626;
  wire seg_18_4_local_g0_1_72344;
  wire seg_18_4_local_g0_2_72345;
  wire seg_18_4_local_g0_3_72346;
  wire seg_18_4_local_g0_4_72347;
  wire seg_18_4_local_g0_6_72349;
  wire seg_18_4_local_g0_7_72350;
  wire seg_18_4_local_g1_0_72351;
  wire seg_18_4_local_g1_1_72352;
  wire seg_18_4_local_g1_2_72353;
  wire seg_18_4_local_g1_3_72354;
  wire seg_18_4_local_g1_4_72355;
  wire seg_18_4_local_g1_5_72356;
  wire seg_18_4_local_g1_7_72358;
  wire seg_18_4_local_g2_0_72359;
  wire seg_18_4_local_g2_1_72360;
  wire seg_18_4_local_g2_5_72364;
  wire seg_18_4_neigh_op_bnl_1_64518;
  wire seg_18_4_neigh_op_bot_0_68348;
  wire seg_18_4_neigh_op_bot_1_68349;
  wire seg_18_4_neigh_op_bot_2_68350;
  wire seg_18_4_neigh_op_bot_3_68351;
  wire seg_18_4_neigh_op_bot_4_68352;
  wire seg_18_4_neigh_op_bot_7_68355;
  wire seg_18_4_neigh_op_tnl_5_64768;
  wire seg_18_4_neigh_op_top_2_68596;
  wire seg_18_4_neigh_op_top_4_68598;
  wire seg_18_4_neigh_op_top_6_68600;
  wire seg_18_4_neigh_op_top_7_68601;
  wire seg_18_4_sp4_h_r_11_72440;
  wire seg_18_4_sp4_h_r_1_72438;
  wire seg_18_4_sp4_h_r_2_72441;
  wire seg_18_4_sp4_h_r_7_72446;
  wire seg_18_4_sp4_r_v_b_45_72458;
  wire seg_18_4_sp4_r_v_b_47_72460;
  wire seg_18_4_sp4_v_b_24_68496;
  wire seg_18_4_sp4_v_b_36_68618;
  wire seg_18_4_sp4_v_b_38_68620;
  wire seg_18_4_sp4_v_b_40_68622;
  wire seg_18_4_sp4_v_b_42_68624;
  wire seg_18_4_sp4_v_b_5_68248;
  wire seg_18_5_glb_netwk_0_5;
  wire seg_18_5_glb_netwk_4_9;
  wire seg_18_5_local_g0_3_72469;
  wire seg_18_5_local_g0_4_72470;
  wire seg_18_5_local_g0_6_72472;
  wire seg_18_5_local_g1_0_72474;
  wire seg_18_5_local_g1_1_72475;
  wire seg_18_5_local_g1_3_72477;
  wire seg_18_5_local_g1_4_72478;
  wire seg_18_5_local_g1_5_72479;
  wire seg_18_5_local_g2_0_72482;
  wire seg_18_5_local_g3_5_72495;
  wire seg_18_5_lutff_2_out_68596;
  wire seg_18_5_lutff_3_out_68597;
  wire seg_18_5_lutff_4_out_68598;
  wire seg_18_5_lutff_5_out_68599;
  wire seg_18_5_lutff_6_out_68600;
  wire seg_18_5_lutff_7_out_68601;
  wire seg_18_5_neigh_op_top_5_68722;
  wire seg_18_5_neigh_op_top_6_68723;
  wire seg_18_5_sp4_h_r_0_72560;
  wire seg_18_5_sp4_h_r_19_68737;
  wire seg_18_5_sp4_h_r_1_72561;
  wire seg_18_5_sp4_h_r_2_72564;
  wire seg_18_5_sp4_h_r_4_72566;
  wire seg_18_5_sp4_h_r_5_72567;
  wire seg_18_5_sp4_h_r_9_72571;
  wire seg_18_5_sp4_r_v_b_8_72212;
  wire seg_18_5_sp4_v_b_16_68499;
  wire seg_18_5_sp4_v_b_20_68503;
  wire seg_18_6_glb_netwk_0_5;
  wire seg_18_6_glb_netwk_4_9;
  wire seg_18_6_local_g0_1_72590;
  wire seg_18_6_local_g0_5_72594;
  wire seg_18_6_local_g1_0_72597;
  wire seg_18_6_local_g1_1_72598;
  wire seg_18_6_local_g1_2_72599;
  wire seg_18_6_local_g1_7_72604;
  wire seg_18_6_local_g2_7_72612;
  wire seg_18_6_local_g3_5_72618;
  wire seg_18_6_lutff_1_out_68718;
  wire seg_18_6_lutff_3_out_68720;
  wire seg_18_6_lutff_5_out_68722;
  wire seg_18_6_lutff_6_out_68723;
  wire seg_18_6_lutff_7_out_68724;
  wire seg_18_6_neigh_op_bnl_5_64768;
  wire seg_18_6_neigh_op_bot_2_68596;
  wire seg_18_6_sp4_h_l_39_57364;
  wire seg_18_6_sp4_h_l_45_57370;
  wire seg_18_6_sp4_h_r_17_68858;
  wire seg_18_6_sp4_h_r_1_72684;
  wire seg_18_6_sp4_h_r_5_72690;
  wire seg_18_6_sp4_h_r_7_72692;
  wire seg_18_6_sp4_h_r_8_72693;
  wire seg_18_6_sp4_r_v_b_15_72452;
  wire seg_18_6_sp4_v_b_0_68496;
  wire seg_18_6_sp4_v_b_21_68627;
  wire seg_18_6_sp4_v_b_31_68747;
  wire seg_18_6_sp4_v_b_8_68504;
  wire seg_18_7_glb_netwk_0_5;
  wire seg_18_7_glb_netwk_4_9;
  wire seg_18_7_local_g0_5_72717;
  wire seg_18_7_local_g0_6_72718;
  wire seg_18_7_local_g0_7_72719;
  wire seg_18_7_local_g1_1_72721;
  wire seg_18_7_local_g1_3_72723;
  wire seg_18_7_local_g1_5_72725;
  wire seg_18_7_local_g1_7_72727;
  wire seg_18_7_local_g2_0_72728;
  wire seg_18_7_local_g2_2_72730;
  wire seg_18_7_local_g2_6_72734;
  wire seg_18_7_local_g3_6_72742;
  wire seg_18_7_neigh_op_bot_7_68724;
  wire seg_18_7_sp12_h_r_14_45988;
  wire seg_18_7_sp12_h_r_16_42156;
  wire seg_18_7_sp12_h_r_18_38326;
  wire seg_18_7_sp12_v_b_18_72435;
  wire seg_18_7_sp4_h_l_43_57491;
  wire seg_18_7_sp4_h_r_11_72809;
  wire seg_18_7_sp4_h_r_14_68980;
  wire seg_18_7_sp4_h_r_20_68986;
  wire seg_18_7_sp4_h_r_28_65150;
  wire seg_18_7_sp4_h_r_2_72810;
  wire seg_18_7_sp4_h_r_3_72811;
  wire seg_18_7_sp4_h_r_40_61320;
  wire seg_18_7_sp4_h_r_42_61322;
  wire seg_18_7_sp4_h_r_46_61316;
  wire seg_18_7_sp4_h_r_6_72814;
  wire seg_18_7_sp4_r_v_b_10_72460;
  wire seg_18_7_sp4_r_v_b_8_72458;
  wire seg_18_7_sp4_v_b_14_68743;
  wire seg_18_7_sp4_v_b_1_68618;
  wire seg_18_7_sp4_v_b_21_68750;
  wire seg_18_7_sp4_v_b_24_68865;
  wire seg_18_7_sp4_v_b_28_68869;
  wire seg_18_7_sp4_v_b_34_68875;
  wire seg_18_7_sp4_v_b_36_68987;
  wire seg_18_7_sp4_v_b_38_68989;
  wire seg_18_7_sp4_v_b_3_68620;
  wire seg_18_7_sp4_v_b_42_68993;
  wire seg_18_7_sp4_v_b_44_68995;
  wire seg_18_7_sp4_v_b_46_68997;
  wire seg_18_7_sp4_v_b_5_68622;
  wire seg_18_7_sp4_v_b_7_68624;
  wire seg_18_7_sp4_v_t_43_69117;
  wire seg_18_8_glb_netwk_0_5;
  wire seg_18_8_glb_netwk_4_9;
  wire seg_18_8_local_g0_1_72836;
  wire seg_18_8_local_g0_5_72840;
  wire seg_18_8_local_g1_3_72846;
  wire seg_18_8_local_g1_5_72848;
  wire seg_18_8_local_g1_7_72850;
  wire seg_18_8_local_g2_3_72854;
  wire seg_18_8_sp4_h_r_0_72929;
  wire seg_18_8_sp4_h_r_18_69107;
  wire seg_18_8_sp4_h_r_21_69108;
  wire seg_18_8_sp4_h_r_2_72933;
  wire seg_18_8_sp4_h_r_32_65277;
  wire seg_18_8_sp4_h_r_40_61443;
  wire seg_18_8_sp4_h_r_46_61439;
  wire seg_18_8_sp4_h_r_5_72936;
  wire seg_18_8_sp4_h_r_9_72940;
  wire seg_18_8_sp4_r_v_b_19_72702;
  wire seg_18_8_sp4_v_b_10_68752;
  wire seg_18_8_sp4_v_b_15_68867;
  wire seg_18_8_sp4_v_b_19_68871;
  wire seg_18_8_sp4_v_b_32_68996;
  wire seg_18_8_sp4_v_b_35_68997;
  wire seg_18_8_sp4_v_b_3_68743;
  wire seg_18_8_sp4_v_t_46_69243;
  wire seg_18_9_glb_netwk_0_5;
  wire seg_18_9_glb_netwk_4_9;
  wire seg_18_9_local_g1_4_72970;
  wire seg_18_9_local_g1_5_72971;
  wire seg_18_9_local_g1_7_72973;
  wire seg_18_9_local_g2_0_72974;
  wire seg_18_9_local_g2_2_72976;
  wire seg_18_9_local_g3_5_72987;
  wire seg_18_9_lutff_0_out_69086;
  wire seg_18_9_lutff_5_out_69091;
  wire seg_18_9_lutff_6_out_69092;
  wire seg_18_9_neigh_op_tnl_2_65380;
  wire seg_18_9_neigh_op_top_4_69213;
  wire seg_18_9_sp4_h_l_42_57738;
  wire seg_18_9_sp4_h_l_46_57732;
  wire seg_18_9_sp4_h_r_15_69225;
  wire seg_18_9_sp4_h_r_34_65392;
  wire seg_18_9_sp4_r_v_b_23_72829;
  wire seg_18_9_sp4_v_b_0_68865;
  wire seg_18_9_sp4_v_b_10_68875;
  wire seg_18_9_sp4_v_b_13_68988;
  wire seg_18_9_sp4_v_b_4_68869;
  wire seg_19_0_local_g1_0_75715;
  wire seg_19_0_local_g1_0_75715_i1;
  wire seg_19_0_local_g1_0_75715_i2;
  wire seg_19_0_local_g1_0_75715_i3;
  wire seg_19_0_span4_horz_r_12_64262;
  wire seg_19_0_span4_vert_0_72044;
  wire seg_19_0_span4_vert_12_72048;
  wire seg_19_10_sp4_v_b_10_72829;
  wire seg_19_10_sp4_v_t_46_73320;
  wire seg_19_11_sp4_h_l_43_61813;
  wire seg_19_11_sp4_v_b_8_72950;
  wire seg_19_12_sp4_h_l_36_61929;
  wire seg_19_12_sp4_h_l_38_61933;
  wire seg_19_12_sp4_h_l_40_61935;
  wire seg_19_12_sp4_h_l_42_61937;
  wire seg_19_12_sp4_h_l_46_61931;
  wire seg_19_17_sp4_h_l_38_62548;
  wire seg_19_1_sp4_h_l_37_60539;
  wire seg_19_1_sp4_h_r_5_75848;
  wire seg_19_2_sp4_h_l_43_60706;
  wire seg_19_2_sp4_h_r_5_75986;
  wire seg_19_2_sp4_v_b_1_72048;
  wire seg_19_3_sp4_h_r_2_76085;
  wire seg_19_4_sp4_h_l_43_60952;
  wire seg_19_5_sp4_h_r_3_76290;
  wire seg_19_5_sp4_h_r_5_76292;
  wire seg_19_6_sp4_h_l_40_61197;
  wire seg_19_6_sp4_h_l_41_61196;
  wire seg_19_6_sp4_h_l_42_61199;
  wire seg_19_7_sp4_h_l_38_61318;
  wire seg_19_7_sp4_h_l_41_61319;
  wire seg_19_7_sp4_v_b_2_72452;
  wire seg_19_8_sp4_h_r_1_76592;
  wire seg_19_9_sp4_v_b_6_72702;
  wire seg_1_10_glb_netwk_0_5;
  wire seg_1_10_glb_netwk_4_9;
  wire seg_1_10_local_g0_3_8081;
  wire seg_1_10_local_g0_5_8083;
  wire seg_1_10_local_g0_7_8085;
  wire seg_1_10_local_g1_3_8089;
  wire seg_1_10_local_g2_1_8095;
  wire seg_1_10_local_g2_4_8098;
  wire seg_1_10_local_g3_2_8104;
  wire seg_1_10_local_g3_6_8108;
  wire seg_1_10_lutff_0_out_1965;
  wire seg_1_10_lutff_1_out_1966;
  wire seg_1_10_lutff_3_out_1968;
  wire seg_1_10_lutff_4_out_1969;
  wire seg_1_10_lutff_5_out_1970;
  wire seg_1_10_lutff_6_out_1971;
  wire seg_1_10_lutff_7_out_1972;
  wire seg_1_10_neigh_op_tnr_1_8185;
  wire seg_1_10_neigh_op_tnr_2_8186;
  wire seg_1_10_neigh_op_tnr_6_8190;
  wire seg_1_10_sp4_h_l_40_2273;
  wire seg_1_10_sp4_h_r_11_8199;
  wire seg_1_10_sp4_h_r_12_2239;
  wire seg_1_10_sp4_h_r_2_8200;
  wire seg_1_10_sp4_h_r_4_8202;
  wire seg_1_10_sp4_h_r_9_8207;
  wire seg_1_10_sp4_r_v_b_13_7915;
  wire seg_1_10_sp4_r_v_b_29_8065;
  wire seg_1_10_sp4_r_v_b_5_7771;
  wire seg_1_10_sp4_v_b_11_1650;
  wire seg_1_10_sp4_v_b_3_1642;
  wire seg_1_10_sp4_v_b_6_1647;
  wire seg_1_10_sp4_v_t_36_2492;
  wire seg_1_10_sp4_v_t_42_2498;
  wire seg_1_10_sp4_v_t_43_2499;
  wire seg_1_10_sp4_v_t_45_2501;
  wire seg_1_11_glb_netwk_0_5;
  wire seg_1_11_glb_netwk_4_9;
  wire seg_1_11_local_g0_3_8228;
  wire seg_1_11_local_g0_7_8232;
  wire seg_1_11_local_g1_2_8235;
  wire seg_1_11_local_g2_5_8246;
  wire seg_1_11_local_g2_6_8247;
  wire seg_1_11_local_g2_7_8248;
  wire seg_1_11_local_g3_3_8252;
  wire seg_1_11_local_g3_5_8254;
  wire seg_1_11_lutff_0_out_2190;
  wire seg_1_11_lutff_1_out_2191;
  wire seg_1_11_lutff_2_out_2192;
  wire seg_1_11_lutff_4_out_2194;
  wire seg_1_11_lutff_5_out_2195;
  wire seg_1_11_lutff_7_out_2197;
  wire seg_1_11_neigh_op_rgt_3_8187;
  wire seg_1_11_sp4_h_l_46_2485;
  wire seg_1_11_sp4_h_r_45_2470;
  wire seg_1_11_sp4_h_r_6_8351;
  wire seg_1_11_sp4_h_r_9_8354;
  wire seg_1_11_sp4_r_v_b_14_8063;
  wire seg_1_11_sp4_r_v_b_23_8072;
  wire seg_1_11_sp4_r_v_b_27_8210;
  wire seg_1_11_sp4_r_v_b_7_7920;
  wire seg_1_11_sp4_v_b_10_1860;
  wire seg_1_11_sp4_v_b_28_2291;
  wire seg_1_11_sp4_v_b_37_2493;
  wire seg_1_11_sp4_v_b_3_1851;
  wire seg_1_11_sp4_v_b_47_2503;
  wire seg_1_11_sp4_v_b_5_1853;
  wire seg_1_11_sp4_v_b_6_1856;
  wire seg_1_11_sp4_v_t_38_2702;
  wire seg_1_11_sp4_v_t_39_2703;
  wire seg_1_12_glb_netwk_0_5;
  wire seg_1_12_glb_netwk_4_9;
  wire seg_1_12_local_g0_3_8375;
  wire seg_1_12_local_g0_5_8377;
  wire seg_1_12_local_g0_6_8378;
  wire seg_1_12_local_g1_0_8380;
  wire seg_1_12_local_g1_3_8383;
  wire seg_1_12_local_g1_4_8384;
  wire seg_1_12_local_g2_4_8392;
  wire seg_1_12_lutff_3_out_2399;
  wire seg_1_12_lutff_5_out_2401;
  wire seg_1_12_lutff_6_out_2402;
  wire seg_1_12_sp4_h_l_38_2684;
  wire seg_1_12_sp4_h_r_12_2653;
  wire seg_1_12_sp4_h_r_19_2696;
  wire seg_1_12_sp4_h_r_24_2657;
  wire seg_1_12_sp4_h_r_36_2670;
  wire seg_1_12_sp4_h_r_4_8496;
  wire seg_1_12_sp4_h_r_5_8497;
  wire seg_1_12_sp4_h_r_6_8498;
  wire seg_1_12_sp4_h_r_8_8500;
  wire seg_1_12_sp4_h_r_9_8501;
  wire seg_1_12_sp4_r_v_b_31_8361;
  wire seg_1_12_sp4_r_v_b_33_8363;
  wire seg_1_12_sp4_v_b_16_2290;
  wire seg_1_12_sp4_v_b_1_2076;
  wire seg_1_12_sp4_v_b_28_2497;
  wire seg_1_12_sp4_v_b_3_2078;
  wire seg_1_12_sp4_v_t_40_2913;
  wire seg_1_13_glb_netwk_0_5;
  wire seg_1_13_glb_netwk_4_9;
  wire seg_1_13_local_g0_0_8519;
  wire seg_1_13_local_g0_3_8522;
  wire seg_1_13_local_g0_6_8525;
  wire seg_1_13_local_g1_0_8527;
  wire seg_1_13_local_g1_2_8529;
  wire seg_1_13_local_g1_4_8531;
  wire seg_1_13_local_g1_6_8533;
  wire seg_1_13_local_g2_0_8535;
  wire seg_1_13_sp4_h_l_38_2893;
  wire seg_1_13_sp4_h_r_0_8637;
  wire seg_1_13_sp4_h_r_1_8638;
  wire seg_1_13_sp4_h_r_22_2864;
  wire seg_1_13_sp4_h_r_26_2868;
  wire seg_1_13_sp4_h_r_28_2870;
  wire seg_1_13_sp4_h_r_2_8641;
  wire seg_1_13_sp4_h_r_30_2872;
  wire seg_1_13_sp4_h_r_4_8643;
  wire seg_1_13_sp4_h_r_5_8644;
  wire seg_1_13_sp4_h_r_8_8647;
  wire seg_1_13_sp4_r_v_b_4_8213;
  wire seg_1_13_sp4_r_v_b_8_8217;
  wire seg_1_13_sp4_v_b_0_2287;
  wire seg_1_13_sp4_v_b_10_2297;
  wire seg_1_13_sp4_v_b_11_2296;
  wire seg_1_13_sp4_v_b_16_2496;
  wire seg_1_13_sp4_v_b_1_2286;
  wire seg_1_13_sp4_v_b_22_2502;
  wire seg_1_13_sp4_v_b_2_2289;
  wire seg_1_13_sp4_v_b_4_2291;
  wire seg_1_13_sp4_v_b_6_2293;
  wire seg_1_13_sp4_v_b_7_2292;
  wire seg_1_13_sp4_v_b_8_2295;
  wire seg_1_13_sp4_v_b_9_2294;
  wire seg_1_13_sp4_v_t_39_3139;
  wire seg_1_14_glb_netwk_0_5;
  wire seg_1_14_glb_netwk_4_9;
  wire seg_1_14_local_g0_3_8669;
  wire seg_1_14_local_g0_4_8670;
  wire seg_1_14_local_g0_5_8671;
  wire seg_1_14_local_g0_7_8673;
  wire seg_1_14_local_g1_6_8680;
  wire seg_1_14_local_g2_1_8683;
  wire seg_1_14_local_g2_2_8684;
  wire seg_1_14_local_g2_7_8689;
  wire seg_1_14_lutff_1_out_2814;
  wire seg_1_14_lutff_3_out_2816;
  wire seg_1_14_lutff_4_out_2817;
  wire seg_1_14_lutff_6_out_2819;
  wire seg_1_14_neigh_op_top_3_3028;
  wire seg_1_14_neigh_op_top_5_3030;
  wire seg_1_14_neigh_op_top_7_3032;
  wire seg_1_14_sp4_h_r_22_3091;
  wire seg_1_14_sp4_h_r_7_8793;
  wire seg_1_14_sp4_r_v_b_15_8505;
  wire seg_1_14_sp4_v_b_0_2493;
  wire seg_1_14_sp4_v_b_10_2503;
  wire seg_1_14_sp4_v_b_26_2912;
  wire seg_1_14_sp4_v_b_2_2495;
  wire seg_1_14_sp4_v_b_31_2915;
  wire seg_1_14_sp4_v_b_33_2917;
  wire seg_1_14_sp4_v_b_3_2494;
  wire seg_1_14_sp4_v_b_4_2497;
  wire seg_1_14_sp4_v_t_38_3348;
  wire seg_1_15_glb_netwk_0_5;
  wire seg_1_15_glb_netwk_4_9;
  wire seg_1_15_local_g0_0_8813;
  wire seg_1_15_local_g1_3_8824;
  wire seg_1_15_local_g1_6_8827;
  wire seg_1_15_local_g2_0_8829;
  wire seg_1_15_local_g2_1_8830;
  wire seg_1_15_local_g2_6_8835;
  wire seg_1_15_local_g3_1_8838;
  wire seg_1_15_local_g3_4_8841;
  wire seg_1_15_lutff_0_out_3025;
  wire seg_1_15_lutff_1_out_3026;
  wire seg_1_15_lutff_2_out_3027;
  wire seg_1_15_lutff_3_out_3028;
  wire seg_1_15_lutff_4_out_3029;
  wire seg_1_15_lutff_5_out_3030;
  wire seg_1_15_lutff_6_out_3031;
  wire seg_1_15_lutff_7_out_3032;
  wire seg_1_15_sp4_h_r_11_8934;
  wire seg_1_15_sp4_v_b_11_2710;
  wire seg_1_15_sp4_v_b_24_3137;
  wire seg_1_15_sp4_v_b_41_3351;
  wire seg_1_15_sp4_v_b_46_3356;
  wire seg_1_15_sp4_v_b_6_2707;
  wire seg_1_15_sp4_v_b_8_2709;
  wire seg_1_15_sp4_v_t_40_3556;
  wire seg_1_15_sp4_v_t_43_3559;
  wire seg_1_15_sp4_v_t_46_3562;
  wire seg_1_16_glb_netwk_0_5;
  wire seg_1_16_glb_netwk_4_9;
  wire seg_1_16_local_g0_5_8965;
  wire seg_1_16_local_g2_1_8977;
  wire seg_1_16_local_g2_5_8981;
  wire seg_1_16_local_g2_6_8982;
  wire seg_1_16_local_g3_0_8984;
  wire seg_1_16_local_g3_4_8988;
  wire seg_1_16_local_g3_5_8989;
  wire seg_1_16_lutff_0_out_3250;
  wire seg_1_16_lutff_2_out_3252;
  wire seg_1_16_lutff_3_out_3253;
  wire seg_1_16_lutff_4_out_3254;
  wire seg_1_16_lutff_5_out_3255;
  wire seg_1_16_lutff_6_out_3256;
  wire seg_1_16_sp4_h_r_2_9082;
  wire seg_1_16_sp4_h_r_8_9088;
  wire seg_1_16_sp4_v_b_10_2920;
  wire seg_1_16_sp4_v_b_29_3350;
  wire seg_1_16_sp4_v_b_33_3354;
  wire seg_1_16_sp4_v_b_37_3553;
  wire seg_1_16_sp4_v_t_36_3760;
  wire seg_1_16_sp4_v_t_39_3763;
  wire seg_1_16_sp4_v_t_41_3765;
  wire seg_1_17_glb_netwk_0_5;
  wire seg_1_17_glb_netwk_4_9;
  wire seg_1_17_local_g0_0_9107;
  wire seg_1_17_local_g0_1_9108;
  wire seg_1_17_local_g0_4_9111;
  wire seg_1_17_local_g2_7_9130;
  wire seg_1_17_lutff_1_out_3457;
  wire seg_1_17_lutff_2_out_3458;
  wire seg_1_17_neigh_op_top_0_3664;
  wire seg_1_17_neigh_op_top_1_3665;
  wire seg_1_17_neigh_op_top_4_3668;
  wire seg_1_17_sp12_v_b_1_7459;
  wire seg_1_17_sp12_v_b_7_7901;
  wire seg_1_17_sp4_h_r_0_9225;
  wire seg_1_17_sp4_r_v_b_7_8802;
  wire seg_1_17_sp4_v_b_14_3348;
  wire seg_1_17_sp4_v_b_47_3771;
  wire seg_1_17_sp4_v_b_4_3141;
  wire seg_1_17_sp4_v_b_5_3140;
  wire seg_1_18_glb_netwk_0_5;
  wire seg_1_18_glb_netwk_4_9;
  wire seg_1_18_local_g0_2_9256;
  wire seg_1_18_local_g0_7_9261;
  wire seg_1_18_local_g1_5_9267;
  wire seg_1_18_local_g3_3_9281;
  wire seg_1_18_lutff_0_out_3664;
  wire seg_1_18_lutff_1_out_3665;
  wire seg_1_18_lutff_4_out_3668;
  wire seg_1_18_lutff_6_out_3670;
  wire seg_1_18_neigh_op_top_5_3878;
  wire seg_1_18_neigh_op_top_7_3880;
  wire seg_1_18_sp4_h_r_10_9374;
  wire seg_1_18_sp4_h_r_1_9373;
  wire seg_1_18_sp4_h_r_2_9376;
  wire seg_1_18_sp4_h_r_8_9382;
  wire seg_1_18_sp4_v_b_2_3349;
  wire seg_1_18_sp4_v_b_43_3976;
  wire seg_1_18_sp4_v_t_40_4200;
  wire seg_1_18_sp4_v_t_46_4206;
  wire seg_1_19_glb_netwk_0_5;
  wire seg_1_19_glb_netwk_4_9;
  wire seg_1_19_local_g0_1_9402;
  wire seg_1_19_local_g0_6_9407;
  wire seg_1_19_local_g1_7_9416;
  wire seg_1_19_lutff_0_out_3873;
  wire seg_1_19_lutff_5_out_3878;
  wire seg_1_19_lutff_7_out_3880;
  wire seg_1_19_neigh_op_top_1_4086;
  wire seg_1_19_neigh_op_top_6_4091;
  wire seg_1_19_neigh_op_top_7_4092;
  wire seg_1_19_sp4_v_t_38_4425;
  wire seg_1_19_sp4_v_t_40_4427;
  wire seg_1_19_sp4_v_t_42_4429;
  wire seg_1_19_sp4_v_t_44_4431;
  wire seg_1_19_sp4_v_t_45_4432;
  wire seg_1_19_sp4_v_t_46_4433;
  wire seg_1_1_glb_netwk_0_5;
  wire seg_1_1_glb_netwk_4_9;
  wire seg_1_1_local_g0_2_6717;
  wire seg_1_1_local_g0_5_6720;
  wire seg_1_1_local_g0_6_6721;
  wire seg_1_1_local_g1_3_6726;
  wire seg_1_1_local_g1_4_6727;
  wire seg_1_1_local_g1_7_6730;
  wire seg_1_1_local_g3_6_6745;
  wire seg_1_1_lutff_2_out_103;
  wire seg_1_1_lutff_5_out_106;
  wire seg_1_1_lutff_6_out_107;
  wire seg_1_1_lutff_7_out_108;
  wire seg_1_1_neigh_op_top_3_119;
  wire seg_1_1_neigh_op_top_6_122;
  wire seg_1_1_sp4_h_r_20_250;
  wire seg_1_1_sp4_r_v_b_29_6871;
  wire seg_1_1_sp4_r_v_b_45_6889;
  wire seg_1_1_sp4_v_b_46_292;
  wire seg_1_20_glb_netwk_0_5;
  wire seg_1_20_glb_netwk_4_9;
  wire seg_1_20_local_g0_6_9554;
  wire seg_1_20_local_g1_4_9560;
  wire seg_1_20_local_g2_0_9564;
  wire seg_1_20_local_g3_4_9576;
  wire seg_1_20_lutff_1_out_4086;
  wire seg_1_20_lutff_2_out_4087;
  wire seg_1_20_lutff_6_out_4091;
  wire seg_1_20_lutff_7_out_4092;
  wire seg_1_20_sp4_v_b_12_3969;
  wire seg_1_20_sp4_v_b_22_3979;
  wire seg_1_20_sp4_v_b_24_4197;
  wire seg_1_20_sp4_v_b_36_4423;
  wire seg_1_20_sp4_v_t_36_4650;
  wire seg_1_20_sp4_v_t_39_4653;
  wire seg_1_20_sp4_v_t_40_4654;
  wire seg_1_20_sp4_v_t_42_4656;
  wire seg_1_20_sp4_v_t_44_4658;
  wire seg_1_20_sp4_v_t_46_4660;
  wire seg_1_21_glb_netwk_0_5;
  wire seg_1_21_glb_netwk_4_9;
  wire seg_1_21_local_g0_5_9700;
  wire seg_1_21_local_g3_2_9721;
  wire seg_1_21_lutff_0_out_4312;
  wire seg_1_21_neigh_op_top_5_4544;
  wire seg_1_21_sp4_h_r_0_9813;
  wire seg_1_21_sp4_h_r_10_9815;
  wire seg_1_21_sp4_h_r_8_9823;
  wire seg_1_21_sp4_v_b_0_3970;
  wire seg_1_21_sp4_v_b_34_4434;
  wire seg_1_21_sp4_v_b_4_3974;
  wire seg_1_21_sp4_v_b_6_3976;
  wire seg_1_21_sp4_v_b_8_3978;
  wire seg_1_21_sp4_v_t_38_4879;
  wire seg_1_21_sp4_v_t_39_4880;
  wire seg_1_21_sp4_v_t_40_4881;
  wire seg_1_22_glb_netwk_0_5;
  wire seg_1_22_glb_netwk_4_9;
  wire seg_1_22_local_g0_1_9843;
  wire seg_1_22_local_g0_6_9848;
  wire seg_1_22_local_g1_1_9851;
  wire seg_1_22_lutff_1_out_4540;
  wire seg_1_22_lutff_5_out_4544;
  wire seg_1_22_sp12_h_r_2_4792;
  wire seg_1_22_sp4_h_r_14_4852;
  wire seg_1_22_sp4_h_r_2_9964;
  wire seg_1_22_sp4_h_r_9_9971;
  wire seg_1_22_sp4_v_b_10_4207;
  wire seg_1_22_sp4_v_b_12_4423;
  wire seg_1_22_sp4_v_b_2_4199;
  wire seg_1_22_sp4_v_b_7_4202;
  wire seg_1_22_sp4_v_b_8_4205;
  wire seg_1_22_sp4_v_t_37_5088;
  wire seg_1_22_sp4_v_t_40_5091;
  wire seg_1_22_sp4_v_t_44_5095;
  wire seg_1_22_sp4_v_t_46_5097;
  wire seg_1_23_glb_netwk_0_5;
  wire seg_1_23_glb_netwk_4_9;
  wire seg_1_23_local_g3_2_10015;
  wire seg_1_23_lutff_2_out_4768;
  wire seg_1_23_sp4_v_b_42_5093;
  wire seg_1_23_sp4_v_t_41_5298;
  wire seg_1_23_sp4_v_t_42_5299;
  wire seg_1_23_sp4_v_t_45_5302;
  wire seg_1_24_sp4_v_t_46_5511;
  wire seg_1_2_glb_netwk_0_5;
  wire seg_1_2_glb_netwk_4_9;
  wire seg_1_2_local_g0_2_6904;
  wire seg_1_2_local_g0_3_6905;
  wire seg_1_2_local_g0_5_6907;
  wire seg_1_2_local_g0_7_6909;
  wire seg_1_2_local_g1_2_6912;
  wire seg_1_2_local_g1_5_6915;
  wire seg_1_2_local_g1_7_6917;
  wire seg_1_2_local_g2_1_6919;
  wire seg_1_2_local_g2_4_6922;
  wire seg_1_2_local_g2_6_6924;
  wire seg_1_2_local_g2_7_6925;
  wire seg_1_2_lutff_1_out_117;
  wire seg_1_2_lutff_2_out_118;
  wire seg_1_2_lutff_3_out_119;
  wire seg_1_2_lutff_4_out_120;
  wire seg_1_2_lutff_5_out_121;
  wire seg_1_2_lutff_6_out_122;
  wire seg_1_2_lutff_7_out_123;
  wire seg_1_2_neigh_op_bot_2_103;
  wire seg_1_2_neigh_op_bot_5_106;
  wire seg_1_2_neigh_op_rgt_1_6826;
  wire seg_1_2_neigh_op_rgt_6_6831;
  wire seg_1_2_neigh_op_rgt_7_6832;
  wire seg_1_2_neigh_op_top_2_453;
  wire seg_1_2_neigh_op_top_5_456;
  wire seg_1_2_neigh_op_top_7_458;
  wire seg_1_2_sp4_h_r_28_523;
  wire seg_1_2_sp4_r_v_b_31_6886;
  wire seg_1_3_glb_netwk_0_5;
  wire seg_1_3_glb_netwk_4_9;
  wire seg_1_3_local_g0_1_7050;
  wire seg_1_3_local_g0_3_7052;
  wire seg_1_3_local_g0_7_7056;
  wire seg_1_3_local_g1_0_7057;
  wire seg_1_3_local_g1_1_7058;
  wire seg_1_3_local_g1_3_7060;
  wire seg_1_3_local_g1_5_7062;
  wire seg_1_3_local_g2_0_7065;
  wire seg_1_3_local_g2_1_7066;
  wire seg_1_3_local_g2_7_7072;
  wire seg_1_3_local_g3_1_7074;
  wire seg_1_3_local_g3_2_7075;
  wire seg_1_3_local_g3_4_7077;
  wire seg_1_3_local_g3_5_7078;
  wire seg_1_3_lutff_0_out_451;
  wire seg_1_3_lutff_1_out_452;
  wire seg_1_3_lutff_2_out_453;
  wire seg_1_3_lutff_3_out_454;
  wire seg_1_3_lutff_4_out_455;
  wire seg_1_3_lutff_5_out_456;
  wire seg_1_3_lutff_6_out_457;
  wire seg_1_3_lutff_7_out_458;
  wire seg_1_3_neigh_op_bnr_0_6825;
  wire seg_1_3_neigh_op_bot_5_121;
  wire seg_1_3_neigh_op_tnr_1_7156;
  wire seg_1_3_neigh_op_top_1_679;
  wire seg_1_3_neigh_op_top_3_681;
  wire seg_1_3_sp4_h_r_10_7169;
  wire seg_1_3_sp4_h_r_20_788;
  wire seg_1_3_sp4_h_r_23_743;
  wire seg_1_3_sp4_h_r_38_761;
  wire seg_1_3_sp4_h_r_8_7177;
  wire seg_1_3_sp4_r_v_b_21_6889;
  wire seg_1_3_sp4_v_b_25_562;
  wire seg_1_4_glb_netwk_0_5;
  wire seg_1_4_glb_netwk_4_9;
  wire seg_1_4_local_g0_0_7196;
  wire seg_1_4_local_g0_3_7199;
  wire seg_1_4_local_g0_5_7201;
  wire seg_1_4_local_g1_1_7205;
  wire seg_1_4_local_g1_3_7207;
  wire seg_1_4_local_g1_5_7209;
  wire seg_1_4_local_g2_1_7213;
  wire seg_1_4_local_g2_2_7214;
  wire seg_1_4_local_g2_6_7218;
  wire seg_1_4_local_g3_2_7222;
  wire seg_1_4_local_g3_6_7226;
  wire seg_1_4_lutff_1_out_679;
  wire seg_1_4_lutff_2_out_680;
  wire seg_1_4_lutff_3_out_681;
  wire seg_1_4_lutff_4_out_682;
  wire seg_1_4_lutff_5_out_683;
  wire seg_1_4_lutff_6_out_684;
  wire seg_1_4_lutff_7_out_685;
  wire seg_1_4_neigh_op_bot_0_451;
  wire seg_1_4_neigh_op_bot_1_452;
  wire seg_1_4_neigh_op_bot_3_454;
  wire seg_1_4_neigh_op_rgt_1_7156;
  wire seg_1_4_neigh_op_rgt_2_7157;
  wire seg_1_4_neigh_op_rgt_6_7161;
  wire seg_1_4_neigh_op_tnr_2_7304;
  wire seg_1_4_neigh_op_top_5_910;
  wire seg_1_4_sp4_v_b_11_292;
  wire seg_1_4_sp4_v_t_37_1227;
  wire seg_1_5_glb_netwk_0_5;
  wire seg_1_5_glb_netwk_4_9;
  wire seg_1_5_local_g0_0_7343;
  wire seg_1_5_local_g0_3_7346;
  wire seg_1_5_local_g0_6_7349;
  wire seg_1_5_local_g1_2_7353;
  wire seg_1_5_local_g1_6_7357;
  wire seg_1_5_local_g2_0_7359;
  wire seg_1_5_local_g2_2_7361;
  wire seg_1_5_local_g2_4_7363;
  wire seg_1_5_local_g2_5_7364;
  wire seg_1_5_local_g2_7_7366;
  wire seg_1_5_lutff_0_out_905;
  wire seg_1_5_lutff_5_out_910;
  wire seg_1_5_lutff_6_out_911;
  wire seg_1_5_neigh_op_bot_6_684;
  wire seg_1_5_neigh_op_rgt_4_7306;
  wire seg_1_5_neigh_op_rgt_7_7309;
  wire seg_1_5_sp4_h_l_38_1210;
  wire seg_1_5_sp4_h_r_10_7463;
  wire seg_1_5_sp4_h_r_14_1201;
  wire seg_1_5_sp4_h_r_18_1223;
  wire seg_1_5_sp4_h_r_20_1225;
  wire seg_1_5_sp4_h_r_22_1181;
  wire seg_1_5_sp4_h_r_3_7466;
  wire seg_1_5_sp4_h_r_4_7467;
  wire seg_1_5_sp4_h_r_6_7469;
  wire seg_1_5_sp4_h_r_8_7471;
  wire seg_1_5_sp4_r_v_b_1_7032;
  wire seg_1_5_sp4_v_b_24_1017;
  wire seg_1_5_sp4_v_b_34_1027;
  wire seg_1_5_sp4_v_b_42_1232;
  wire seg_1_5_sp4_v_b_46_1236;
  wire seg_1_5_sp4_v_b_8_571;
  wire seg_1_5_sp4_v_t_38_1434;
  wire seg_1_6_glb_netwk_0_5;
  wire seg_1_6_glb_netwk_4_9;
  wire seg_1_6_local_g0_1_7491;
  wire seg_1_6_local_g2_0_7506;
  wire seg_1_6_local_g2_3_7509;
  wire seg_1_6_local_g2_4_7510;
  wire seg_1_6_local_g3_5_7519;
  wire seg_1_6_lutff_1_out_1131;
  wire seg_1_6_lutff_3_out_1133;
  wire seg_1_6_lutff_5_out_1135;
  wire seg_1_6_lutff_6_out_1136;
  wire seg_1_6_neigh_op_rgt_0_7449;
  wire seg_1_6_neigh_op_rgt_3_7452;
  wire seg_1_6_neigh_op_rgt_4_7453;
  wire seg_1_6_sp12_v_b_22_7459;
  wire seg_1_6_sp4_h_l_44_1423;
  wire seg_1_6_sp4_h_r_2_7612;
  wire seg_1_6_sp4_h_r_7_7617;
  wire seg_1_6_sp4_h_r_9_7619;
  wire seg_1_6_sp4_v_b_40_1436;
  wire seg_1_6_sp4_v_b_44_1440;
  wire seg_1_6_sp4_v_b_8_798;
  wire seg_1_6_sp4_v_t_41_1645;
  wire seg_1_7_glb_netwk_0_5;
  wire seg_1_7_local_g1_3_7648;
  wire seg_1_7_local_g1_6_7651;
  wire seg_1_7_lutff_1_out_1337;
  wire seg_1_7_sp4_h_r_10_7757;
  wire seg_1_7_sp4_h_r_11_7758;
  wire seg_1_7_sp4_h_r_2_7759;
  wire seg_1_7_sp4_h_r_6_7763;
  wire seg_1_7_sp4_v_b_0_1017;
  wire seg_1_7_sp4_v_b_10_1027;
  wire seg_1_7_sp4_v_b_2_1019;
  wire seg_1_7_sp4_v_b_6_1023;
  wire seg_1_7_sp4_v_t_43_1856;
  wire seg_1_7_sp4_v_t_44_1857;
  wire seg_1_8_glb_netwk_0_5;
  wire seg_1_8_glb_netwk_4_9;
  wire seg_1_8_local_g1_0_7792;
  wire seg_1_8_local_g1_6_7798;
  wire seg_1_8_local_g2_1_7801;
  wire seg_1_8_local_g2_2_7802;
  wire seg_1_8_local_g2_6_7806;
  wire seg_1_8_local_g3_0_7808;
  wire seg_1_8_local_g3_4_7812;
  wire seg_1_8_local_g3_7_7815;
  wire seg_1_8_lutff_0_out_1544;
  wire seg_1_8_lutff_1_out_1545;
  wire seg_1_8_lutff_2_out_1546;
  wire seg_1_8_lutff_3_out_1547;
  wire seg_1_8_lutff_4_out_1548;
  wire seg_1_8_lutff_6_out_1550;
  wire seg_1_8_lutff_7_out_1551;
  wire seg_1_8_sp12_h_r_0_7898;
  wire seg_1_8_sp4_h_r_10_7904;
  wire seg_1_8_sp4_h_r_28_1810;
  wire seg_1_8_sp4_h_r_5_7909;
  wire seg_1_8_sp4_v_b_16_1436;
  wire seg_1_8_sp4_v_b_30_1647;
  wire seg_1_8_sp4_v_b_38_1851;
  wire seg_1_8_sp4_v_b_39_1852;
  wire seg_1_8_sp4_v_b_3_1228;
  wire seg_1_8_sp4_v_b_40_1853;
  wire seg_1_8_sp4_v_b_46_1859;
  wire seg_1_8_sp4_v_b_6_1233;
  wire seg_1_8_sp4_v_b_8_1235;
  wire seg_1_8_sp4_v_t_46_2086;
  wire seg_1_9_glb_netwk_0_5;
  wire seg_1_9_glb_netwk_4_9;
  wire seg_1_9_local_g0_0_7931;
  wire seg_1_9_local_g0_5_7936;
  wire seg_1_9_local_g1_5_7944;
  wire seg_1_9_local_g1_7_7946;
  wire seg_1_9_local_g3_1_7956;
  wire seg_1_9_local_g3_5_7960;
  wire seg_1_9_local_g3_6_7961;
  wire seg_1_9_local_g3_7_7962;
  wire seg_1_9_lutff_5_out_1758;
  wire seg_1_9_lutff_7_out_1760;
  wire seg_1_9_neigh_op_top_0_1965;
  wire seg_1_9_sp12_h_r_13_1992;
  wire seg_1_9_sp12_h_r_5_2002;
  wire seg_1_9_sp4_h_r_16_2071;
  wire seg_1_9_sp4_h_r_25_2032;
  wire seg_1_9_sp4_h_r_4_8055;
  wire seg_1_9_sp4_h_r_6_8057;
  wire seg_1_9_sp4_h_r_8_8059;
  wire seg_1_9_sp4_r_v_b_22_7777;
  wire seg_1_9_sp4_r_v_b_23_7778;
  wire seg_1_9_sp4_r_v_b_29_7918;
  wire seg_1_9_sp4_r_v_b_41_8066;
  wire seg_1_9_sp4_r_v_b_45_8070;
  wire seg_1_9_sp4_v_b_10_1443;
  wire seg_1_9_sp4_v_b_11_1442;
  wire seg_1_9_sp4_v_b_15_1643;
  wire seg_1_9_sp4_v_b_24_1850;
  wire seg_1_9_sp4_v_b_32_1858;
  wire seg_1_9_sp4_v_b_34_1860;
  wire seg_1_9_sp4_v_b_36_2076;
  wire seg_1_9_sp4_v_b_38_2078;
  wire seg_1_9_sp4_v_b_45_2085;
  wire seg_1_9_sp4_v_b_8_1441;
  wire seg_1_9_sp4_v_b_9_1440;
  wire seg_1_9_sp4_v_t_38_2288;
  wire seg_1_9_sp4_v_t_41_2291;
  wire seg_20_10_glb_netwk_0_5;
  wire seg_20_10_glb_netwk_4_9;
  wire seg_20_10_local_g0_1_80113;
  wire seg_20_10_local_g0_2_80114;
  wire seg_20_10_local_g0_6_80118;
  wire seg_20_10_local_g0_7_80119;
  wire seg_20_10_local_g1_6_80126;
  wire seg_20_10_local_g1_7_80127;
  wire seg_20_10_lutff_0_out_76651;
  wire seg_20_10_lutff_1_out_76652;
  wire seg_20_10_lutff_5_out_76656;
  wire seg_20_10_neigh_op_bot_7_76556;
  wire seg_20_10_neigh_op_top_6_76759;
  wire seg_20_10_sp4_h_l_39_65517;
  wire seg_20_10_sp4_h_l_40_65520;
  wire seg_20_10_sp4_h_l_43_65521;
  wire seg_20_10_sp4_h_r_1_80207;
  wire seg_20_10_sp4_h_r_23_76797;
  wire seg_20_10_sp4_h_r_24_73175;
  wire seg_20_10_sp4_h_r_26_73179;
  wire seg_20_10_sp4_h_r_6_80214;
  wire seg_20_10_sp4_h_r_8_80216;
  wire seg_20_10_sp4_v_b_11_76511;
  wire seg_20_10_sp4_v_b_18_76609;
  wire seg_20_11_glb_netwk_0_5;
  wire seg_20_11_glb_netwk_4_9;
  wire seg_20_11_local_g0_7_80242;
  wire seg_20_11_local_g1_1_80244;
  wire seg_20_11_lutff_6_out_76759;
  wire seg_20_11_neigh_op_bot_1_76652;
  wire seg_20_11_sp4_h_r_15_76901;
  wire seg_20_11_sp4_h_r_30_73306;
  wire seg_20_12_glb_netwk_0_5;
  wire seg_20_12_glb_netwk_1_6;
  wire seg_20_12_glb_netwk_4_9;
  wire seg_20_12_local_g0_4_80362;
  wire seg_20_12_local_g3_1_80383;
  wire seg_20_12_sp4_h_r_20_77010;
  wire seg_20_12_sp4_v_b_25_76909;
  wire seg_20_12_sp4_v_b_4_76710;
  wire seg_20_14_glb_netwk_0_5;
  wire seg_20_14_local_g1_3_80615;
  wire seg_20_14_local_g3_3_80631;
  wire seg_20_14_sp4_h_l_42_66014;
  wire seg_20_14_sp4_h_r_38_69841;
  wire seg_20_14_sp4_r_v_b_19_80471;
  wire seg_20_14_sp4_v_b_19_77018;
  wire seg_20_15_sp4_h_l_37_66128;
  wire seg_20_2_glb_netwk_0_5;
  wire seg_20_2_glb_netwk_4_9;
  wire seg_20_2_local_g0_2_79130;
  wire seg_20_2_local_g1_7_79143;
  wire seg_20_2_local_g3_3_79155;
  wire seg_20_2_lutff_2_out_75801;
  wire seg_20_2_lutff_7_out_75806;
  wire seg_20_2_sp4_h_l_38_64534;
  wire seg_20_2_sp4_h_l_47_64531;
  wire seg_20_2_sp4_h_r_36_68361;
  wire seg_20_2_sp4_h_r_46_68363;
  wire seg_20_2_sp4_v_b_27_75885;
  wire seg_20_3_glb_netwk_0_5;
  wire seg_20_3_glb_netwk_4_9;
  wire seg_20_3_local_g1_0_79259;
  wire seg_20_3_local_g1_1_79260;
  wire seg_20_3_local_g2_1_79268;
  wire seg_20_3_local_g2_3_79270;
  wire seg_20_3_local_g3_3_79278;
  wire seg_20_3_local_g3_4_79279;
  wire seg_20_3_lutff_0_out_75937;
  wire seg_20_3_lutff_1_out_75938;
  wire seg_20_3_neigh_op_rgt_3_79213;
  wire seg_20_3_sp4_h_l_41_64658;
  wire seg_20_3_sp4_h_l_43_64660;
  wire seg_20_3_sp4_h_r_28_72320;
  wire seg_20_3_sp4_h_r_38_68488;
  wire seg_20_3_sp4_h_r_42_68492;
  wire seg_20_3_sp4_h_r_46_68486;
  wire seg_20_3_sp4_h_r_4_79351;
  wire seg_20_3_sp4_r_v_b_11_79104;
  wire seg_20_3_sp4_r_v_b_20_79114;
  wire seg_20_3_sp4_r_v_b_25_79234;
  wire seg_20_4_glb_netwk_0_5;
  wire seg_20_4_glb_netwk_4_9;
  wire seg_20_4_local_g1_5_79387;
  wire seg_20_4_local_g1_6_79388;
  wire seg_20_4_local_g3_3_79401;
  wire seg_20_4_sp4_h_l_38_64780;
  wire seg_20_4_sp4_h_r_18_76192;
  wire seg_20_4_sp4_h_r_5_79475;
  wire seg_20_4_sp4_h_r_6_79476;
  wire seg_20_4_sp4_h_r_7_79477;
  wire seg_20_4_sp4_r_v_b_19_79241;
  wire seg_20_4_sp4_v_b_13_75992;
  wire seg_20_4_sp4_v_b_43_76202;
  wire seg_20_5_glb_netwk_0_5;
  wire seg_20_5_glb_netwk_4_9;
  wire seg_20_5_local_g0_4_79501;
  wire seg_20_5_local_g0_7_79504;
  wire seg_20_5_local_g1_0_79505;
  wire seg_20_5_local_g1_3_79508;
  wire seg_20_5_local_g2_6_79519;
  wire seg_20_5_local_g3_1_79522;
  wire seg_20_5_local_g3_6_79527;
  wire seg_20_5_local_g3_7_79528;
  wire seg_20_5_sp4_h_l_43_64906;
  wire seg_20_5_sp4_h_l_45_64908;
  wire seg_20_5_sp4_h_r_16_76292;
  wire seg_20_5_sp4_h_r_28_72566;
  wire seg_20_5_sp4_h_r_2_79595;
  wire seg_20_5_sp4_h_r_36_68730;
  wire seg_20_5_sp4_h_r_38_68734;
  wire seg_20_5_sp4_h_r_40_68736;
  wire seg_20_5_sp4_h_r_42_68738;
  wire seg_20_5_sp4_h_r_46_68732;
  wire seg_20_5_sp4_h_r_5_79598;
  wire seg_20_5_sp4_h_r_8_79601;
  wire seg_20_5_sp4_r_v_b_14_79359;
  wire seg_20_5_sp4_r_v_b_22_79367;
  wire seg_20_5_sp4_r_v_b_23_79368;
  wire seg_20_5_sp4_r_v_b_27_79482;
  wire seg_20_5_sp4_r_v_b_41_79608;
  wire seg_20_5_sp4_v_b_12_76093;
  wire seg_20_5_sp4_v_b_15_76096;
  wire seg_20_5_sp4_v_t_41_76404;
  wire seg_20_6_glb_netwk_0_5;
  wire seg_20_6_glb_netwk_4_9;
  wire seg_20_6_local_g1_2_79630;
  wire seg_20_6_local_g1_3_79631;
  wire seg_20_6_local_g1_4_79632;
  wire seg_20_6_local_g1_5_79633;
  wire seg_20_6_local_g2_4_79640;
  wire seg_20_6_local_g2_5_79641;
  wire seg_20_6_local_g2_6_79642;
  wire seg_20_6_local_g3_1_79645;
  wire seg_20_6_local_g3_2_79646;
  wire seg_20_6_local_g3_3_79647;
  wire seg_20_6_local_g3_5_79649;
  wire seg_20_6_sp4_h_l_40_65028;
  wire seg_20_6_sp4_h_l_41_65027;
  wire seg_20_6_sp4_h_l_43_65029;
  wire seg_20_6_sp4_h_l_45_65031;
  wire seg_20_6_sp4_h_r_18_76396;
  wire seg_20_6_sp4_h_r_1_79715;
  wire seg_20_6_sp4_h_r_2_79718;
  wire seg_20_6_sp4_h_r_32_72693;
  wire seg_20_6_sp4_h_r_34_72685;
  wire seg_20_6_sp4_h_r_37_68852;
  wire seg_20_6_sp4_h_r_3_79719;
  wire seg_20_6_sp4_h_r_40_68859;
  wire seg_20_6_sp4_h_r_43_68860;
  wire seg_20_6_sp4_h_r_45_68862;
  wire seg_20_6_sp4_r_v_b_5_79361;
  wire seg_20_6_sp4_v_b_12_76195;
  wire seg_20_6_sp4_v_b_26_76300;
  wire seg_20_6_sp4_v_b_33_76305;
  wire seg_20_6_sp4_v_b_36_76399;
  wire seg_20_6_sp4_v_b_3_76095;
  wire seg_20_6_sp4_v_b_46_76409;
  wire seg_20_6_sp4_v_t_41_76506;
  wire seg_20_7_glb_netwk_0_5;
  wire seg_20_7_glb_netwk_4_9;
  wire seg_20_7_local_g0_2_79745;
  wire seg_20_7_local_g0_7_79750;
  wire seg_20_7_local_g1_1_79752;
  wire seg_20_7_local_g1_6_79757;
  wire seg_20_7_local_g3_3_79770;
  wire seg_20_7_sp4_h_l_38_65149;
  wire seg_20_7_sp4_h_l_40_65151;
  wire seg_20_7_sp4_h_l_42_65153;
  wire seg_20_7_sp4_h_l_43_65152;
  wire seg_20_7_sp4_h_l_45_65154;
  wire seg_20_7_sp4_h_l_47_65146;
  wire seg_20_7_sp4_h_r_42_68984;
  wire seg_20_7_sp4_h_r_7_79846;
  wire seg_20_7_sp4_h_r_9_79848;
  wire seg_20_7_sp4_r_v_b_43_79856;
  wire seg_20_7_sp4_v_b_10_76206;
  wire seg_20_7_sp4_v_b_11_76205;
  wire seg_20_7_sp4_v_b_22_76307;
  wire seg_20_8_glb_netwk_0_5;
  wire seg_20_8_glb_netwk_4_9;
  wire seg_20_8_local_g3_3_79893;
  wire seg_20_8_neigh_op_tnr_3_79951;
  wire seg_20_8_sp4_h_l_38_65272;
  wire seg_20_8_sp4_h_l_46_65270;
  wire seg_20_8_sp4_h_r_12_76592;
  wire seg_20_8_sp4_v_b_28_76506;
  wire seg_20_8_sp4_v_b_2_76300;
  wire seg_20_8_sp4_v_t_41_76710;
  wire seg_20_9_glb_netwk_0_5;
  wire seg_20_9_glb_netwk_4_9;
  wire seg_20_9_local_g0_7_79996;
  wire seg_20_9_local_g1_1_79998;
  wire seg_20_9_local_g1_7_80004;
  wire seg_20_9_local_g3_7_80020;
  wire seg_20_9_lutff_7_out_76556;
  wire seg_20_9_neigh_op_bnr_1_79826;
  wire seg_20_9_neigh_op_bnr_7_79832;
  wire seg_20_9_neigh_op_rgt_7_79955;
  wire seg_20_9_sp4_h_l_47_65392;
  wire seg_20_9_sp4_h_r_42_69230;
  wire seg_20_9_sp4_h_r_8_80093;
  wire seg_20_9_sp4_h_r_9_80094;
  wire seg_20_9_sp4_v_b_15_76504;
  wire seg_20_9_sp4_v_b_22_76511;
  wire seg_21_0_local_g1_4_82750;
  wire seg_21_0_span4_vert_36_79105;
  wire seg_21_10_glb_netwk_0_5;
  wire seg_21_10_glb_netwk_4_9;
  wire seg_21_10_local_g0_0_83943;
  wire seg_21_10_local_g1_0_83951;
  wire seg_21_10_local_g1_3_83954;
  wire seg_21_10_local_g1_5_83956;
  wire seg_21_10_local_g1_7_83958;
  wire seg_21_10_lutff_2_out_80073;
  wire seg_21_10_lutff_3_out_80074;
  wire seg_21_10_neigh_op_bot_0_79948;
  wire seg_21_10_neigh_op_lft_0_76651;
  wire seg_21_10_neigh_op_lft_5_76656;
  wire seg_21_10_sp4_h_l_36_69345;
  wire seg_21_10_sp4_h_l_38_69349;
  wire seg_21_10_sp4_h_l_42_69353;
  wire seg_21_10_sp4_h_l_44_69355;
  wire seg_21_10_sp4_h_l_46_69347;
  wire seg_21_10_sp4_h_r_0_84037;
  wire seg_21_10_sp4_h_r_2_84041;
  wire seg_21_10_sp4_h_r_40_73182;
  wire seg_21_10_sp4_h_r_5_84044;
  wire seg_21_10_sp4_v_b_15_79975;
  wire seg_21_10_sp4_v_b_19_79979;
  wire seg_21_10_sp4_v_b_2_79852;
  wire seg_21_10_sp4_v_b_7_79855;
  wire seg_21_11_sp4_h_l_41_69473;
  wire seg_21_11_sp4_h_l_45_69477;
  wire seg_21_11_sp4_h_l_47_69469;
  wire seg_21_11_sp4_h_r_2_84164;
  wire seg_21_11_sp4_v_b_3_79974;
  wire seg_21_12_sp4_h_l_38_69595;
  wire seg_21_12_sp4_h_l_40_69597;
  wire seg_21_12_sp4_h_l_42_69599;
  wire seg_21_13_sp4_h_l_37_69713;
  wire seg_21_13_sp4_h_l_40_69720;
  wire seg_21_13_sp4_h_l_41_69719;
  wire seg_21_13_sp4_h_l_45_69723;
  wire seg_21_13_sp4_h_l_47_69715;
  wire seg_21_2_sp4_h_l_37_68360;
  wire seg_21_3_glb_netwk_0_5;
  wire seg_21_3_glb_netwk_4_9;
  wire seg_21_3_local_g2_2_83100;
  wire seg_21_3_local_g2_4_83102;
  wire seg_21_3_local_g3_0_83106;
  wire seg_21_3_local_g3_6_83112;
  wire seg_21_3_lutff_3_out_79213;
  wire seg_21_3_neigh_op_rgt_0_83041;
  wire seg_21_3_neigh_op_rgt_2_83043;
  wire seg_21_3_neigh_op_tnr_6_83170;
  wire seg_21_3_sp4_h_l_36_68484;
  wire seg_21_3_sp4_h_r_0_83176;
  wire seg_21_3_sp4_h_r_2_83180;
  wire seg_21_3_sp4_h_r_36_72315;
  wire seg_21_3_sp4_h_r_46_72317;
  wire seg_21_3_sp4_h_r_6_83184;
  wire seg_21_3_sp4_r_v_b_12_82936;
  wire seg_21_4_glb_netwk_0_5;
  wire seg_21_4_glb_netwk_4_9;
  wire seg_21_4_local_g0_1_83206;
  wire seg_21_4_local_g1_6_83219;
  wire seg_21_4_local_g2_6_83227;
  wire seg_21_4_local_g2_7_83228;
  wire seg_21_4_local_g3_7_83236;
  wire seg_21_4_neigh_op_rgt_7_83171;
  wire seg_21_4_neigh_op_tnr_6_83293;
  wire seg_21_4_sp4_h_l_36_68607;
  wire seg_21_4_sp4_h_l_37_68606;
  wire seg_21_4_sp4_h_l_39_68610;
  wire seg_21_4_sp4_h_l_43_68614;
  wire seg_21_4_sp4_h_r_16_79475;
  wire seg_21_4_sp4_h_r_18_79477;
  wire seg_21_4_sp4_h_r_1_83300;
  wire seg_21_4_sp4_h_r_36_72438;
  wire seg_21_4_sp4_h_r_3_83304;
  wire seg_21_4_sp4_h_r_42_72446;
  wire seg_21_4_sp4_h_r_46_72440;
  wire seg_21_4_sp4_h_r_4_83305;
  wire seg_21_4_sp4_h_r_6_83307;
  wire seg_21_4_sp4_v_b_39_79483;
  wire seg_21_5_glb_netwk_0_5;
  wire seg_21_5_glb_netwk_4_9;
  wire seg_21_5_local_g0_0_83328;
  wire seg_21_5_local_g3_4_83356;
  wire seg_21_5_local_g3_5_83357;
  wire seg_21_5_neigh_op_rgt_4_83291;
  wire seg_21_5_sp4_h_l_37_68729;
  wire seg_21_5_sp4_h_l_39_68733;
  wire seg_21_5_sp4_h_l_44_68740;
  wire seg_21_5_sp4_h_r_1_83423;
  wire seg_21_5_sp4_h_r_36_72561;
  wire seg_21_5_sp4_h_r_3_83427;
  wire seg_21_5_sp4_h_r_40_72567;
  wire seg_21_5_sp4_h_r_44_72571;
  wire seg_21_5_sp4_r_v_b_24_83312;
  wire seg_21_5_sp4_v_b_45_79612;
  wire seg_21_5_sp4_v_b_6_79241;
  wire seg_21_6_glb_netwk_0_5;
  wire seg_21_6_glb_netwk_4_9;
  wire seg_21_6_local_g0_1_83452;
  wire seg_21_6_local_g2_4_83471;
  wire seg_21_6_local_g3_4_83479;
  wire seg_21_6_local_g3_6_83481;
  wire seg_21_6_lutff_6_out_79585;
  wire seg_21_6_neigh_op_rgt_4_83414;
  wire seg_21_6_sp4_h_l_36_68853;
  wire seg_21_6_sp4_h_r_10_83547;
  wire seg_21_6_sp4_h_r_14_79719;
  wire seg_21_6_sp4_h_r_1_83546;
  wire seg_21_6_sp4_h_r_3_83550;
  wire seg_21_6_sp4_h_r_40_72690;
  wire seg_21_6_sp4_h_r_42_72692;
  wire seg_21_6_sp4_h_r_6_83553;
  wire seg_21_6_sp4_r_v_b_25_83434;
  wire seg_21_6_sp4_v_b_36_79726;
  wire seg_21_7_glb_netwk_0_5;
  wire seg_21_7_glb_netwk_4_9;
  wire seg_21_7_local_g0_2_83576;
  wire seg_21_7_local_g0_3_83577;
  wire seg_21_7_local_g0_5_83579;
  wire seg_21_7_local_g3_2_83600;
  wire seg_21_7_lutff_1_out_79703;
  wire seg_21_7_lutff_2_out_79704;
  wire seg_21_7_neigh_op_tnr_2_83658;
  wire seg_21_7_sp4_h_l_38_68980;
  wire seg_21_7_sp4_h_r_0_83668;
  wire seg_21_7_sp4_h_r_10_83670;
  wire seg_21_7_sp4_h_r_2_83672;
  wire seg_21_7_sp4_h_r_38_72811;
  wire seg_21_7_sp4_h_r_3_83673;
  wire seg_21_7_sp4_h_r_46_72809;
  wire seg_21_7_sp4_r_v_b_33_83565;
  wire seg_21_7_sp4_v_b_13_79604;
  wire seg_21_8_glb_netwk_0_5;
  wire seg_21_8_glb_netwk_4_9;
  wire seg_21_8_local_g0_2_83699;
  wire seg_21_8_local_g0_4_83701;
  wire seg_21_8_local_g0_6_83703;
  wire seg_21_8_local_g0_7_83704;
  wire seg_21_8_local_g1_1_83706;
  wire seg_21_8_local_g1_2_83707;
  wire seg_21_8_local_g1_5_83710;
  wire seg_21_8_local_g1_6_83711;
  wire seg_21_8_local_g2_3_83716;
  wire seg_21_8_local_g2_4_83717;
  wire seg_21_8_local_g2_6_83719;
  wire seg_21_8_local_g2_7_83720;
  wire seg_21_8_local_g3_0_83721;
  wire seg_21_8_local_g3_4_83725;
  wire seg_21_8_local_g3_5_83726;
  wire seg_21_8_local_g3_6_83727;
  wire seg_21_8_lutff_1_out_79826;
  wire seg_21_8_lutff_7_out_79832;
  wire seg_21_8_neigh_op_bnr_2_83535;
  wire seg_21_8_neigh_op_bnr_4_83537;
  wire seg_21_8_neigh_op_bnr_5_83538;
  wire seg_21_8_neigh_op_bnr_7_83540;
  wire seg_21_8_neigh_op_bot_1_79703;
  wire seg_21_8_neigh_op_bot_2_79704;
  wire seg_21_8_neigh_op_rgt_0_83656;
  wire seg_21_8_neigh_op_rgt_3_83659;
  wire seg_21_8_neigh_op_rgt_4_83660;
  wire seg_21_8_neigh_op_rgt_5_83661;
  wire seg_21_8_neigh_op_rgt_6_83662;
  wire seg_21_8_neigh_op_tnr_4_83783;
  wire seg_21_8_neigh_op_tnr_6_83785;
  wire seg_21_8_neigh_op_tnr_7_83786;
  wire seg_21_8_neigh_op_top_6_79954;
  wire seg_21_8_sp12_h_r_12_61432;
  wire seg_21_8_sp12_h_r_14_57603;
  wire seg_21_8_sp4_h_r_0_83791;
  wire seg_21_8_sp4_h_r_40_72936;
  wire seg_21_8_sp4_h_r_44_72940;
  wire seg_21_8_sp4_h_r_4_83797;
  wire seg_21_8_sp4_h_r_5_83798;
  wire seg_21_8_sp4_h_r_6_83799;
  wire seg_21_8_sp4_h_r_8_83801;
  wire seg_21_8_sp4_v_b_26_79852;
  wire seg_21_9_glb_netwk_0_5;
  wire seg_21_9_glb_netwk_4_9;
  wire seg_21_9_local_g0_5_83825;
  wire seg_21_9_local_g1_2_83830;
  wire seg_21_9_local_g1_3_83831;
  wire seg_21_9_local_g1_4_83832;
  wire seg_21_9_local_g1_6_83834;
  wire seg_21_9_local_g1_7_83835;
  wire seg_21_9_local_g2_0_83836;
  wire seg_21_9_local_g2_4_83840;
  wire seg_21_9_local_g3_3_83847;
  wire seg_21_9_local_g3_6_83850;
  wire seg_21_9_lutff_0_out_79948;
  wire seg_21_9_lutff_3_out_79951;
  wire seg_21_9_lutff_4_out_79952;
  wire seg_21_9_lutff_6_out_79954;
  wire seg_21_9_lutff_7_out_79955;
  wire seg_21_9_neigh_op_bnr_5_83661;
  wire seg_21_9_neigh_op_rgt_0_83779;
  wire seg_21_9_neigh_op_rgt_3_83782;
  wire seg_21_9_neigh_op_top_2_80073;
  wire seg_21_9_neigh_op_top_3_80074;
  wire seg_21_9_sp4_h_r_14_80088;
  wire seg_21_9_sp4_h_r_20_80094;
  wire seg_21_9_sp4_h_r_3_83919;
  wire seg_21_9_sp4_h_r_5_83921;
  wire seg_21_9_sp4_h_r_8_83924;
  wire seg_21_9_sp4_r_v_b_12_83680;
  wire seg_21_9_sp4_v_b_18_79855;
  wire seg_21_9_sp4_v_b_23_79860;
  wire seg_21_9_sp4_v_b_9_79734;
  wire seg_22_0_local_g1_6_86583;
  wire seg_22_0_span4_vert_22_82921;
  wire seg_22_10_sp12_h_r_18_54019;
  wire seg_22_10_sp4_h_l_39_73179;
  wire seg_22_10_sp4_h_r_11_87871;
  wire seg_22_10_sp4_h_r_1_87869;
  wire seg_22_10_sp4_h_r_32_80216;
  wire seg_22_10_sp4_h_r_3_87873;
  wire seg_22_11_sp4_h_r_11_87994;
  wire seg_22_11_sp4_h_r_1_87992;
  wire seg_22_12_sp4_h_r_11_88117;
  wire seg_22_12_sp4_h_r_5_88121;
  wire seg_22_13_sp4_h_r_3_88242;
  wire seg_22_13_sp4_h_r_5_88244;
  wire seg_22_13_sp4_h_r_9_88248;
  wire seg_22_2_sp4_v_t_46_83198;
  wire seg_22_3_glb_netwk_0_5;
  wire seg_22_3_glb_netwk_4_9;
  wire seg_22_3_local_g0_4_86917;
  wire seg_22_3_local_g1_3_86924;
  wire seg_22_3_local_g3_3_86940;
  wire seg_22_3_lutff_0_out_83041;
  wire seg_22_3_lutff_2_out_83043;
  wire seg_22_3_sp4_h_r_11_87010;
  wire seg_22_3_sp4_h_r_8_87017;
  wire seg_22_3_sp4_v_b_20_82945;
  wire seg_22_3_sp4_v_b_35_83075;
  wire seg_22_3_sp4_v_t_46_83321;
  wire seg_22_4_glb_netwk_0_5;
  wire seg_22_4_glb_netwk_4_9;
  wire seg_22_4_local_g0_0_87036;
  wire seg_22_4_local_g2_2_87054;
  wire seg_22_4_local_g2_7_87059;
  wire seg_22_4_lutff_6_out_83170;
  wire seg_22_4_lutff_7_out_83171;
  wire seg_22_4_neigh_op_tnr_7_87125;
  wire seg_22_4_sp12_h_r_12_64771;
  wire seg_22_4_sp4_h_r_0_87130;
  wire seg_22_4_sp4_v_b_42_83317;
  wire seg_22_4_sp4_v_t_40_83438;
  wire seg_22_4_sp4_v_t_42_83440;
  wire seg_22_4_sp4_v_t_44_83442;
  wire seg_22_5_glb_netwk_0_5;
  wire seg_22_5_glb_netwk_4_9;
  wire seg_22_5_local_g0_4_87163;
  wire seg_22_5_local_g2_1_87176;
  wire seg_22_5_local_g2_2_87177;
  wire seg_22_5_local_g2_3_87178;
  wire seg_22_5_local_g3_0_87183;
  wire seg_22_5_lutff_4_out_83291;
  wire seg_22_5_lutff_6_out_83293;
  wire seg_22_5_neigh_op_rgt_0_87118;
  wire seg_22_5_neigh_op_rgt_1_87119;
  wire seg_22_5_neigh_op_tnr_3_87244;
  wire seg_22_5_sp4_h_r_11_87256;
  wire seg_22_5_sp4_h_r_14_83427;
  wire seg_22_5_sp4_h_r_1_87254;
  wire seg_22_5_sp4_h_r_20_83433;
  wire seg_22_5_sp4_h_r_32_79601;
  wire seg_22_5_sp4_h_r_38_76290;
  wire seg_22_5_sp4_h_r_3_87258;
  wire seg_22_5_sp4_h_r_7_87262;
  wire seg_22_5_sp4_h_r_9_87264;
  wire seg_22_5_sp4_v_b_26_83314;
  wire seg_22_5_sp4_v_t_46_83567;
  wire seg_22_6_glb_netwk_0_5;
  wire seg_22_6_glb_netwk_4_9;
  wire seg_22_6_local_g2_3_87301;
  wire seg_22_6_local_g2_7_87305;
  wire seg_22_6_lutff_4_out_83414;
  wire seg_22_6_neigh_op_rgt_7_87248;
  wire seg_22_6_sp12_h_r_16_57356;
  wire seg_22_6_sp4_h_l_46_72686;
  wire seg_22_6_sp4_h_r_12_83546;
  wire seg_22_6_sp4_h_r_1_87377;
  wire seg_22_6_sp4_h_r_5_87383;
  wire seg_22_6_sp4_v_b_43_83564;
  wire seg_22_6_sp4_v_t_45_83689;
  wire seg_22_7_glb_netwk_0_5;
  wire seg_22_7_glb_netwk_4_9;
  wire seg_22_7_local_g1_0_87413;
  wire seg_22_7_local_g2_7_87428;
  wire seg_22_7_local_g3_1_87430;
  wire seg_22_7_local_g3_5_87434;
  wire seg_22_7_lutff_2_out_83535;
  wire seg_22_7_lutff_4_out_83537;
  wire seg_22_7_lutff_5_out_83538;
  wire seg_22_7_lutff_7_out_83540;
  wire seg_22_7_sp4_h_r_11_87502;
  wire seg_22_7_sp4_h_r_7_87508;
  wire seg_22_7_sp4_h_r_9_87510;
  wire seg_22_7_sp4_r_v_b_24_87389;
  wire seg_22_7_sp4_v_b_25_83557;
  wire seg_22_7_sp4_v_b_29_83561;
  wire seg_22_7_sp4_v_b_31_83563;
  wire seg_22_7_sp4_v_t_41_83808;
  wire seg_22_8_glb_netwk_0_5;
  wire seg_22_8_glb_netwk_4_9;
  wire seg_22_8_local_g1_3_87539;
  wire seg_22_8_local_g1_6_87542;
  wire seg_22_8_local_g1_7_87543;
  wire seg_22_8_local_g2_3_87547;
  wire seg_22_8_local_g2_6_87550;
  wire seg_22_8_local_g3_5_87557;
  wire seg_22_8_lutff_0_out_83656;
  wire seg_22_8_lutff_2_out_83658;
  wire seg_22_8_lutff_3_out_83659;
  wire seg_22_8_lutff_4_out_83660;
  wire seg_22_8_lutff_5_out_83661;
  wire seg_22_8_lutff_6_out_83662;
  wire seg_22_8_sp4_h_r_5_87629;
  wire seg_22_8_sp4_h_r_7_87631;
  wire seg_22_8_sp4_h_r_9_87633;
  wire seg_22_8_sp4_r_v_b_21_87397;
  wire seg_22_8_sp4_r_v_b_27_87513;
  wire seg_22_8_sp4_v_b_14_83559;
  wire seg_22_8_sp4_v_b_15_83560;
  wire seg_22_8_sp4_v_b_30_83687;
  wire seg_22_8_sp4_v_b_35_83690;
  wire seg_22_8_sp4_v_t_40_83930;
  wire seg_22_9_glb_netwk_0_5;
  wire seg_22_9_glb_netwk_4_9;
  wire seg_22_9_local_g1_6_87665;
  wire seg_22_9_local_g2_1_87668;
  wire seg_22_9_local_g3_1_87676;
  wire seg_22_9_local_g3_2_87677;
  wire seg_22_9_local_g3_7_87682;
  wire seg_22_9_lutff_0_out_83779;
  wire seg_22_9_lutff_3_out_83782;
  wire seg_22_9_lutff_4_out_83783;
  wire seg_22_9_lutff_6_out_83785;
  wire seg_22_9_lutff_7_out_83786;
  wire seg_22_9_sp4_r_v_b_17_87516;
  wire seg_22_9_sp4_r_v_b_18_87517;
  wire seg_22_9_sp4_r_v_b_23_87522;
  wire seg_22_9_sp4_v_b_14_83682;
  wire seg_22_9_sp4_v_b_25_83803;
  wire seg_22_9_sp4_v_t_39_84052;
  wire seg_22_9_sp4_v_t_45_84058;
  wire seg_22_9_sp4_v_t_47_84060;
  wire seg_23_0_local_g1_2_90410;
  wire seg_23_0_span4_vert_0_86737;
  wire seg_23_0_span4_vert_16_86745;
  wire seg_23_0_span4_vert_19_86748;
  wire seg_23_0_span4_vert_37_86768;
  wire seg_23_0_span4_vert_42_86774;
  wire seg_23_10_sp4_h_r_0_91699;
  wire seg_23_10_sp4_h_r_10_91701;
  wire seg_23_10_sp4_h_r_2_91703;
  wire seg_23_10_sp4_h_r_4_91705;
  wire seg_23_11_sp4_h_l_43_76905;
  wire seg_23_12_sp4_h_l_40_77006;
  wire seg_23_12_sp4_h_l_42_77008;
  wire seg_23_12_sp4_h_l_43_77007;
  wire seg_23_12_sp4_h_l_46_77002;
  wire seg_23_12_sp4_h_r_4_91951;
  wire seg_23_13_sp4_h_r_6_92076;
  wire seg_23_1_sp4_v_b_0_86737;
  wire seg_23_2_sp4_h_l_43_75987;
  wire seg_23_2_sp4_v_b_5_86745;
  wire seg_23_3_sp4_v_t_39_87145;
  wire seg_23_4_sp4_h_l_42_76192;
  wire seg_23_4_sp4_h_l_43_76191;
  wire seg_23_5_glb_netwk_0_5;
  wire seg_23_5_glb_netwk_4_9;
  wire seg_23_5_local_g0_1_90991;
  wire seg_23_5_local_g2_3_91009;
  wire seg_23_5_local_g3_0_91014;
  wire seg_23_5_local_g3_4_91018;
  wire seg_23_5_local_g3_7_91021;
  wire seg_23_5_lutff_0_out_87118;
  wire seg_23_5_lutff_1_out_87119;
  wire seg_23_5_lutff_7_out_87125;
  wire seg_23_5_neigh_op_top_1_87242;
  wire seg_23_5_sp4_h_r_0_91084;
  wire seg_23_5_sp4_h_r_31_83431;
  wire seg_23_5_sp4_h_r_35_83425;
  wire seg_23_5_sp4_h_r_40_79598;
  wire seg_23_5_sp4_h_r_8_91094;
  wire seg_23_5_sp4_v_b_24_87143;
  wire seg_23_5_sp4_v_b_26_87145;
  wire seg_23_5_sp4_v_b_36_87265;
  wire seg_23_6_glb_netwk_0_5;
  wire seg_23_6_glb_netwk_4_9;
  wire seg_23_6_local_g2_4_91133;
  wire seg_23_6_local_g3_0_91137;
  wire seg_23_6_local_g3_4_91141;
  wire seg_23_6_lutff_1_out_87242;
  wire seg_23_6_lutff_3_out_87244;
  wire seg_23_6_lutff_7_out_87248;
  wire seg_23_6_sp4_h_l_36_76388;
  wire seg_23_6_sp4_h_l_47_76389;
  wire seg_23_6_sp4_h_r_10_91209;
  wire seg_23_6_sp4_h_r_8_91217;
  wire seg_23_6_sp4_r_v_b_40_91223;
  wire seg_23_6_sp4_v_b_28_87270;
  wire seg_23_6_sp4_v_b_44_87396;
  wire seg_23_6_sp4_v_b_6_87026;
  wire seg_23_7_sp4_h_l_42_76498;
  wire seg_23_7_sp4_h_l_43_76497;
  wire seg_23_7_sp4_h_r_0_91330;
  wire seg_23_8_glb_netwk_0_5;
  wire seg_23_8_glb_netwk_4_9;
  wire seg_23_8_local_g2_5_91380;
  wire seg_23_8_sp4_h_r_30_83799;
  wire seg_23_8_sp4_h_r_8_91463;
  wire seg_23_8_sp4_v_b_29_87515;
  wire seg_23_8_sp4_v_t_41_87762;
  wire seg_23_9_glb_netwk_0_5;
  wire seg_23_9_glb_netwk_4_9;
  wire seg_23_9_local_g1_5_91495;
  wire seg_23_9_sp4_h_r_38_80088;
  wire seg_23_9_sp4_v_b_21_87520;
  wire seg_23_9_sp4_v_t_43_87887;
  wire seg_24_0_span4_vert_13_90573;
  wire seg_24_13_sp4_h_r_9_96090;
  wire seg_24_2_sp4_h_l_43_79230;
  wire seg_24_6_sp4_h_l_40_79721;
  wire seg_24_6_sp4_h_l_42_79723;
  wire seg_24_6_sp4_h_l_44_79725;
  wire seg_24_6_sp4_h_l_46_79717;
  wire seg_24_6_sp4_h_r_11_95109;
  wire seg_24_6_sp4_h_r_1_95107;
  wire seg_24_7_sp4_h_l_38_79842;
  wire seg_24_7_sp4_h_l_40_79844;
  wire seg_24_7_sp4_h_l_41_79843;
  wire seg_24_7_sp4_h_l_47_79839;
  wire seg_24_9_sp4_v_t_44_91719;
  wire seg_25_10_sp4_h_l_38_84042;
  wire seg_25_10_sp4_h_l_41_84043;
  wire seg_25_10_sp4_h_l_42_84046;
  wire seg_25_10_sp4_h_l_44_84048;
  wire seg_25_10_sp4_h_l_45_84047;
  wire seg_25_10_sp4_h_l_46_84040;
  wire seg_25_10_sp4_h_l_47_84039;
  wire seg_25_10_sp4_h_r_24_91699;
  wire seg_25_10_sp4_h_r_26_91703;
  wire seg_25_10_sp4_h_r_28_91705;
  wire seg_25_10_sp4_h_r_34_91701;
  wire seg_25_10_sp4_h_r_36_87869;
  wire seg_25_10_sp4_h_r_38_87873;
  wire seg_25_10_sp4_h_r_46_87871;
  wire seg_25_10_sp4_v_b_0_95258;
  wire seg_25_11_local_g0_0_100150;
  wire seg_25_11_local_g0_4_100154;
  wire seg_25_11_local_g0_5_100155;
  wire seg_25_11_local_g0_6_100156;
  wire seg_25_11_local_g1_6_100164;
  wire seg_25_11_local_g2_2_100168;
  wire seg_25_11_local_g2_3_100169;
  wire seg_25_11_local_g2_4_100170;
  wire seg_25_11_local_g2_5_100171;
  wire seg_25_11_local_g2_6_100172;
  wire seg_25_11_local_g2_7_100173;
  wire seg_25_11_local_g3_1_100175;
  wire seg_25_11_local_g3_2_100176;
  wire seg_25_11_local_g3_4_100178;
  wire seg_25_11_local_g3_6_100180;
  wire seg_25_11_local_g3_7_100181;
  wire seg_25_11_sp4_h_l_41_84166;
  wire seg_25_11_sp4_h_l_43_84168;
  wire seg_25_11_sp4_h_l_45_84170;
  wire seg_25_11_sp4_h_r_0_100236;
  wire seg_25_11_sp4_h_r_26_91826;
  wire seg_25_11_sp4_h_r_2_100240;
  wire seg_25_11_sp4_h_r_36_87992;
  wire seg_25_11_sp4_h_r_46_87994;
  wire seg_25_11_sp4_h_r_4_100242;
  wire seg_25_11_sp4_h_r_6_100244;
  wire seg_25_11_sp4_v_b_0_95397;
  wire seg_25_11_sp4_v_b_10_95407;
  wire seg_25_11_sp4_v_b_12_95535;
  wire seg_25_11_sp4_v_b_14_95537;
  wire seg_25_11_sp4_v_b_21_95544;
  wire seg_25_11_sp4_v_b_22_95545;
  wire seg_25_11_sp4_v_b_27_95676;
  wire seg_25_11_sp4_v_b_28_95679;
  wire seg_25_11_sp4_v_b_30_95681;
  wire seg_25_11_sp4_v_b_31_95680;
  wire seg_25_11_sp4_v_b_38_95815;
  wire seg_25_11_sp4_v_b_39_95816;
  wire seg_25_11_sp4_v_b_41_95818;
  wire seg_25_11_sp4_v_b_42_95819;
  wire seg_25_11_sp4_v_b_44_95821;
  wire seg_25_11_sp4_v_b_45_95822;
  wire seg_25_11_sp4_v_b_8_95405;
  wire seg_25_12_local_g0_2_100302;
  wire seg_25_12_local_g0_3_100303;
  wire seg_25_12_local_g1_1_100309;
  wire seg_25_12_local_g1_2_100310;
  wire seg_25_12_local_g1_3_100311;
  wire seg_25_12_local_g1_4_100312;
  wire seg_25_12_local_g1_5_100313;
  wire seg_25_12_local_g1_6_100314;
  wire seg_25_12_local_g2_1_100317;
  wire seg_25_12_local_g2_2_100318;
  wire seg_25_12_local_g2_3_100319;
  wire seg_25_12_local_g2_4_100320;
  wire seg_25_12_local_g3_1_100325;
  wire seg_25_12_local_g3_2_100326;
  wire seg_25_12_local_g3_6_100330;
  wire seg_25_12_local_g3_7_100331;
  wire seg_25_12_sp4_h_l_38_84288;
  wire seg_25_12_sp4_h_l_45_84293;
  wire seg_25_12_sp4_h_l_46_84286;
  wire seg_25_12_sp4_h_r_25_91946;
  wire seg_25_12_sp4_h_r_28_91951;
  wire seg_25_12_sp4_h_r_2_100391;
  wire seg_25_12_sp4_h_r_30_91953;
  wire seg_25_12_sp4_h_r_31_91954;
  wire seg_25_12_sp4_h_r_35_91948;
  wire seg_25_12_sp4_h_r_3_100392;
  wire seg_25_12_sp4_h_r_40_88121;
  wire seg_25_12_sp4_h_r_46_88117;
  wire seg_25_12_sp4_h_r_4_100393;
  wire seg_25_12_sp4_v_b_10_95546;
  wire seg_25_12_sp4_v_b_14_95676;
  wire seg_25_12_sp4_v_b_16_95678;
  wire seg_25_12_sp4_v_b_17_95679;
  wire seg_25_12_sp4_v_b_18_95680;
  wire seg_25_12_sp4_v_b_19_95681;
  wire seg_25_12_sp4_v_b_20_95682;
  wire seg_25_12_sp4_v_b_21_95683;
  wire seg_25_12_sp4_v_b_26_95816;
  wire seg_25_12_sp4_v_b_2_95538;
  wire seg_25_12_sp4_v_b_33_95821;
  wire seg_25_12_sp4_v_b_34_95824;
  wire seg_25_12_sp4_v_b_36_95952;
  wire seg_25_12_sp4_v_b_6_95542;
  wire seg_25_13_sp4_h_l_36_84407;
  wire seg_25_13_sp4_h_l_38_84411;
  wire seg_25_13_sp4_h_l_41_84412;
  wire seg_25_13_sp4_h_l_43_84414;
  wire seg_25_13_sp4_h_l_45_84416;
  wire seg_25_13_sp4_h_r_20_96090;
  wire seg_25_13_sp4_h_r_30_92076;
  wire seg_25_13_sp4_h_r_38_88242;
  wire seg_25_13_sp4_h_r_40_88244;
  wire seg_25_13_sp4_h_r_44_88248;
  wire seg_25_13_sp4_v_b_0_95675;
  wire seg_25_13_sp4_v_b_10_95685;
  wire seg_25_13_sp4_v_b_2_95677;
  wire seg_25_3_sp4_h_l_36_83177;
  wire seg_25_3_sp4_v_b_10_94273;
  wire seg_25_3_sp4_v_t_37_94841;
  wire seg_25_3_sp4_v_t_39_94843;
  wire seg_25_4_sp4_h_l_39_83303;
  wire seg_25_4_sp4_h_l_44_83310;
  wire seg_25_4_sp4_h_l_45_83309;
  wire seg_25_4_sp4_h_l_47_83301;
  wire seg_25_4_sp4_v_b_2_90451;
  wire seg_25_4_sp4_v_b_3_90450;
  wire seg_25_4_sp4_v_t_36_94979;
  wire seg_25_4_sp4_v_t_41_94984;
  wire seg_25_4_sp4_v_t_43_94986;
  wire seg_25_4_sp4_v_t_44_94987;
  wire seg_25_5_sp4_h_l_37_83422;
  wire seg_25_5_sp4_h_l_40_83429;
  wire seg_25_5_sp4_h_l_45_83432;
  wire seg_25_5_sp4_h_r_24_91084;
  wire seg_25_5_sp4_h_r_32_91094;
  wire seg_25_5_sp4_h_r_36_87254;
  wire seg_25_5_sp4_h_r_38_87258;
  wire seg_25_5_sp4_h_r_42_87262;
  wire seg_25_5_sp4_h_r_44_87264;
  wire seg_25_5_sp4_h_r_46_87256;
  wire seg_25_5_sp4_v_b_34_94851;
  wire seg_25_5_sp4_v_t_36_95118;
  wire seg_25_5_sp4_v_t_38_95120;
  wire seg_25_5_sp4_v_t_42_95124;
  wire seg_25_5_sp4_v_t_46_95128;
  wire seg_25_6_local_g0_0_99370;
  wire seg_25_6_local_g0_3_99373;
  wire seg_25_6_local_g1_2_99380;
  wire seg_25_6_local_g1_5_99383;
  wire seg_25_6_local_g1_7_99385;
  wire seg_25_6_local_g2_0_99386;
  wire seg_25_6_local_g2_2_99388;
  wire seg_25_6_local_g2_3_99389;
  wire seg_25_6_local_g2_5_99391;
  wire seg_25_6_local_g3_0_99394;
  wire seg_25_6_local_g3_1_99395;
  wire seg_25_6_local_g3_2_99396;
  wire seg_25_6_local_g3_4_99398;
  wire seg_25_6_local_g3_5_99399;
  wire seg_25_6_local_g3_6_99400;
  wire seg_25_6_local_g3_7_99401;
  wire seg_25_6_sp4_h_l_44_83556;
  wire seg_25_6_sp4_h_r_10_99458;
  wire seg_25_6_sp4_h_r_12_95107;
  wire seg_25_6_sp4_h_r_13_95106;
  wire seg_25_6_sp4_h_r_16_95113;
  wire seg_25_6_sp4_h_r_18_95115;
  wire seg_25_6_sp4_h_r_22_95109;
  wire seg_25_6_sp4_h_r_23_95108;
  wire seg_25_6_sp4_h_r_24_91207;
  wire seg_25_6_sp4_h_r_25_91208;
  wire seg_25_6_sp4_h_r_28_91213;
  wire seg_25_6_sp4_h_r_32_91217;
  wire seg_25_6_sp4_h_r_34_91209;
  wire seg_25_6_sp4_h_r_36_87377;
  wire seg_25_6_sp4_h_r_40_87383;
  wire seg_25_6_sp4_h_r_46_87379;
  wire seg_25_6_sp4_v_b_19_94847;
  wire seg_25_6_sp4_v_b_26_94982;
  wire seg_25_6_sp4_v_b_27_94981;
  wire seg_25_6_sp4_v_b_30_94986;
  wire seg_25_6_sp4_v_b_32_94988;
  wire seg_25_6_sp4_v_b_34_94990;
  wire seg_25_6_sp4_v_b_37_95119;
  wire seg_25_6_sp4_v_b_45_95127;
  wire seg_25_6_sp4_v_b_47_95129;
  wire seg_25_6_sp4_v_t_38_95259;
  wire seg_25_6_sp4_v_t_43_95264;
  wire seg_25_7_local_g0_0_99520;
  wire seg_25_7_local_g0_1_99521;
  wire seg_25_7_local_g0_3_99523;
  wire seg_25_7_local_g0_7_99527;
  wire seg_25_7_local_g1_1_99529;
  wire seg_25_7_local_g1_2_99530;
  wire seg_25_7_local_g1_4_99532;
  wire seg_25_7_local_g1_5_99533;
  wire seg_25_7_local_g1_6_99534;
  wire seg_25_7_local_g1_7_99535;
  wire seg_25_7_local_g2_0_99536;
  wire seg_25_7_local_g2_7_99543;
  wire seg_25_7_local_g3_0_99544;
  wire seg_25_7_local_g3_1_99545;
  wire seg_25_7_local_g3_3_99547;
  wire seg_25_7_local_g3_5_99549;
  wire seg_25_7_sp12_h_r_20_61309;
  wire seg_25_7_sp4_h_r_17_95251;
  wire seg_25_7_sp4_h_r_19_95253;
  wire seg_25_7_sp4_h_r_21_95255;
  wire seg_25_7_sp4_h_r_23_95247;
  wire seg_25_7_sp4_h_r_24_91330;
  wire seg_25_7_sp4_h_r_27_91335;
  wire seg_25_7_sp4_h_r_33_91341;
  wire seg_25_7_sp4_h_r_42_87508;
  wire seg_25_7_sp4_h_r_44_87510;
  wire seg_25_7_sp4_h_r_46_87502;
  wire seg_25_7_sp4_v_b_0_94841;
  wire seg_25_7_sp4_v_b_10_94851;
  wire seg_25_7_sp4_v_b_15_94982;
  wire seg_25_7_sp4_v_b_16_94983;
  wire seg_25_7_sp4_v_b_18_94985;
  wire seg_25_7_sp4_v_b_1_94840;
  wire seg_25_7_sp4_v_b_20_94987;
  wire seg_25_7_sp4_v_b_24_95119;
  wire seg_25_7_sp4_v_b_29_95122;
  wire seg_25_7_sp4_v_b_2_94843;
  wire seg_25_7_sp4_v_b_32_95127;
  wire seg_25_7_sp4_v_b_38_95259;
  wire seg_25_7_sp4_v_b_39_95260;
  wire seg_25_7_sp4_v_b_6_94847;
  wire seg_25_7_sp4_v_t_37_95397;
  wire seg_25_7_sp4_v_t_45_95405;
  wire seg_25_7_sp4_v_t_47_95407;
  wire seg_25_8_sp4_h_r_32_91463;
  wire seg_25_8_sp4_h_r_40_87629;
  wire seg_25_8_sp4_h_r_42_87631;
  wire seg_25_8_sp4_h_r_44_87633;
  wire seg_25_8_sp4_v_b_18_95124;
  wire seg_25_8_sp4_v_b_22_95128;
  wire seg_25_8_sp4_v_b_30_95264;
  wire seg_25_8_sp4_v_b_4_94984;
  wire seg_25_8_sp4_v_t_36_95535;
  wire seg_25_8_sp4_v_t_39_95538;
  wire seg_25_8_sp4_v_t_43_95542;
  wire seg_25_8_sp4_v_t_46_95545;
  wire seg_25_8_sp4_v_t_47_95546;
  wire seg_25_9_sp4_v_t_37_95675;
  wire seg_25_9_sp4_v_t_39_95677;
  wire seg_25_9_sp4_v_t_40_95678;
  wire seg_25_9_sp4_v_t_44_95682;
  wire seg_25_9_sp4_v_t_47_95685;
  wire seg_2_10_glb_netwk_0_5;
  wire seg_2_10_glb_netwk_5_10;
  wire seg_2_10_local_g0_1_12419;
  wire seg_2_10_local_g1_6_12432;
  wire seg_2_10_local_g1_7_12433;
  wire seg_2_10_local_g2_2_12436;
  wire seg_2_10_local_g2_5_12439;
  wire seg_2_10_local_g3_0_12442;
  wire seg_2_10_local_g3_1_12443;
  wire seg_2_10_local_g3_4_12446;
  wire seg_2_10_lutff_0_out_8037;
  wire seg_2_10_lutff_2_out_8039;
  wire seg_2_10_lutff_4_out_8041;
  wire seg_2_10_lutff_6_out_8043;
  wire seg_2_10_lutff_7_out_8044;
  wire seg_2_10_neigh_op_lft_6_1971;
  wire seg_2_10_neigh_op_tnl_0_2190;
  wire seg_2_10_neigh_op_tnl_1_2191;
  wire seg_2_10_neigh_op_tnl_4_2194;
  wire seg_2_10_neigh_op_tnl_5_2195;
  wire seg_2_10_sp4_h_r_10_12514;
  wire seg_2_10_sp4_h_r_11_12515;
  wire seg_2_10_sp4_h_r_1_12513;
  wire seg_2_10_sp4_h_r_2_12516;
  wire seg_2_10_sp4_h_r_42_2248;
  wire seg_2_10_sp4_r_v_b_37_12525;
  wire seg_2_10_sp4_r_v_b_7_12161;
  wire seg_2_10_sp4_v_t_36_8355;
  wire seg_2_10_sp4_v_t_42_8361;
  wire seg_2_10_sp4_v_t_43_8362;
  wire seg_2_10_sp4_v_t_44_8363;
  wire seg_2_10_sp4_v_t_45_8364;
  wire seg_2_11_glb_netwk_0_5;
  wire seg_2_11_glb_netwk_4_9;
  wire seg_2_11_local_g0_0_12541;
  wire seg_2_11_local_g0_1_12542;
  wire seg_2_11_local_g0_3_12544;
  wire seg_2_11_local_g0_5_12546;
  wire seg_2_11_local_g1_4_12553;
  wire seg_2_11_local_g1_5_12554;
  wire seg_2_11_local_g1_7_12556;
  wire seg_2_11_local_g2_2_12559;
  wire seg_2_11_local_g2_6_12563;
  wire seg_2_11_local_g2_7_12564;
  wire seg_2_11_local_g3_0_12565;
  wire seg_2_11_local_g3_1_12566;
  wire seg_2_11_local_g3_2_12567;
  wire seg_2_11_local_g3_3_12568;
  wire seg_2_11_local_g3_4_12569;
  wire seg_2_11_local_g3_5_12570;
  wire seg_2_11_lutff_1_out_8185;
  wire seg_2_11_lutff_2_out_8186;
  wire seg_2_11_lutff_3_out_8187;
  wire seg_2_11_lutff_5_out_8189;
  wire seg_2_11_lutff_6_out_8190;
  wire seg_2_11_neigh_op_bot_4_8041;
  wire seg_2_11_neigh_op_tnr_1_12624;
  wire seg_2_11_neigh_op_tnr_2_12625;
  wire seg_2_11_neigh_op_tnr_3_12626;
  wire seg_2_11_neigh_op_tnr_4_12627;
  wire seg_2_11_neigh_op_tnr_5_12628;
  wire seg_2_11_neigh_op_tnr_6_12629;
  wire seg_2_11_neigh_op_tnr_7_12630;
  wire seg_2_11_sp4_h_r_10_12637;
  wire seg_2_11_sp4_h_r_16_8350;
  wire seg_2_11_sp4_h_r_17_8349;
  wire seg_2_11_sp4_h_r_21_8353;
  wire seg_2_11_sp4_h_r_23_8345;
  wire seg_2_11_sp4_h_r_4_12641;
  wire seg_2_11_sp4_h_r_6_12643;
  wire seg_2_11_sp4_h_r_8_12645;
  wire seg_2_11_sp4_h_r_9_12646;
  wire seg_2_11_sp4_r_v_b_27_12526;
  wire seg_2_11_sp4_r_v_b_29_12528;
  wire seg_2_11_sp4_r_v_b_31_12530;
  wire seg_2_11_sp4_r_v_b_47_12658;
  wire seg_2_11_sp4_v_b_24_8209;
  wire seg_2_11_sp4_v_b_26_8211;
  wire seg_2_11_sp4_v_b_5_7918;
  wire seg_2_11_sp4_v_b_8_7923;
  wire seg_2_11_sp4_v_t_39_8505;
  wire seg_2_12_glb_netwk_0_5;
  wire seg_2_12_glb_netwk_4_9;
  wire seg_2_12_local_g0_3_12667;
  wire seg_2_12_local_g0_5_12669;
  wire seg_2_12_local_g2_1_12681;
  wire seg_2_12_local_g2_3_12683;
  wire seg_2_12_local_g2_5_12685;
  wire seg_2_12_local_g3_0_12688;
  wire seg_2_12_local_g3_2_12690;
  wire seg_2_12_local_g3_4_12692;
  wire seg_2_12_local_g3_7_12695;
  wire seg_2_12_lutff_0_out_8331;
  wire seg_2_12_lutff_1_out_8332;
  wire seg_2_12_lutff_2_out_8333;
  wire seg_2_12_lutff_3_out_8334;
  wire seg_2_12_lutff_4_out_8335;
  wire seg_2_12_lutff_5_out_8336;
  wire seg_2_12_lutff_6_out_8337;
  wire seg_2_12_neigh_op_rgt_7_12630;
  wire seg_2_12_sp4_h_l_36_2670;
  wire seg_2_12_sp4_h_r_11_12761;
  wire seg_2_12_sp4_h_r_27_2675;
  wire seg_2_12_sp4_h_r_29_2695;
  wire seg_2_12_sp4_h_r_32_2698;
  wire seg_2_12_sp4_h_r_33_2699;
  wire seg_2_12_sp4_h_r_3_12763;
  wire seg_2_12_sp4_h_r_6_12766;
  wire seg_2_12_sp4_h_r_8_12768;
  wire seg_2_12_sp4_r_v_b_20_12532;
  wire seg_2_12_sp4_r_v_b_27_12649;
  wire seg_2_12_sp4_r_v_b_29_12651;
  wire seg_2_12_sp4_r_v_b_31_12653;
  wire seg_2_12_sp4_v_b_10_8072;
  wire seg_2_12_sp4_v_b_11_8071;
  wire seg_2_12_sp4_v_b_26_8358;
  wire seg_2_12_sp4_v_b_4_8066;
  wire seg_2_12_sp4_v_b_8_8070;
  wire seg_2_13_glb_netwk_0_5;
  wire seg_2_13_glb_netwk_4_9;
  wire seg_2_13_local_g0_3_12790;
  wire seg_2_13_local_g0_6_12793;
  wire seg_2_13_local_g1_3_12798;
  wire seg_2_13_local_g1_7_12802;
  wire seg_2_13_local_g2_1_12804;
  wire seg_2_13_local_g2_7_12810;
  wire seg_2_13_local_g3_1_12812;
  wire seg_2_13_local_g3_3_12814;
  wire seg_2_13_local_g3_5_12816;
  wire seg_2_13_local_g3_7_12818;
  wire seg_2_13_lutff_0_out_8478;
  wire seg_2_13_lutff_1_out_8479;
  wire seg_2_13_lutff_4_out_8482;
  wire seg_2_13_lutff_6_out_8484;
  wire seg_2_13_lutff_7_out_8485;
  wire seg_2_13_neigh_op_bnr_7_12630;
  wire seg_2_13_neigh_op_tnl_1_2814;
  wire seg_2_13_neigh_op_tnl_3_2816;
  wire seg_2_13_neigh_op_tnr_5_12874;
  wire seg_2_13_sp4_h_l_37_2878;
  wire seg_2_13_sp4_h_r_10_12883;
  wire seg_2_13_sp4_h_r_14_8642;
  wire seg_2_13_sp4_h_r_19_8645;
  wire seg_2_13_sp4_h_r_26_2873;
  wire seg_2_13_sp4_h_r_4_12887;
  wire seg_2_13_sp4_h_r_6_12889;
  wire seg_2_13_sp4_r_v_b_11_12534;
  wire seg_2_13_sp4_r_v_b_23_12658;
  wire seg_2_13_sp4_v_b_10_8219;
  wire seg_2_13_sp4_v_b_11_8218;
  wire seg_2_13_sp4_v_b_12_8355;
  wire seg_2_13_sp4_v_t_42_8802;
  wire seg_2_14_glb_netwk_0_5;
  wire seg_2_14_glb_netwk_4_9;
  wire seg_2_14_local_g0_3_12913;
  wire seg_2_14_local_g1_1_12919;
  wire seg_2_14_local_g1_2_12920;
  wire seg_2_14_local_g1_7_12925;
  wire seg_2_14_local_g2_1_12927;
  wire seg_2_14_local_g2_2_12928;
  wire seg_2_14_local_g2_5_12931;
  wire seg_2_14_local_g2_6_12932;
  wire seg_2_14_local_g3_0_12934;
  wire seg_2_14_local_g3_1_12935;
  wire seg_2_14_neigh_op_bnr_7_12753;
  wire seg_2_14_neigh_op_rgt_0_12869;
  wire seg_2_14_neigh_op_rgt_1_12870;
  wire seg_2_14_neigh_op_top_1_8773;
  wire seg_2_14_neigh_op_top_2_8774;
  wire seg_2_14_neigh_op_top_3_8775;
  wire seg_2_14_sp4_h_r_10_13006;
  wire seg_2_14_sp4_h_r_12_8785;
  wire seg_2_14_sp4_h_r_25_3089;
  wire seg_2_14_sp4_h_r_26_3100;
  wire seg_2_14_sp4_h_r_36_3092;
  wire seg_2_14_sp4_r_v_b_14_12772;
  wire seg_2_14_sp4_r_v_b_31_12899;
  wire seg_2_14_sp4_r_v_b_35_12903;
  wire seg_2_14_sp4_v_b_45_8805;
  wire seg_2_14_sp4_v_b_6_8362;
  wire seg_2_14_sp4_v_b_8_8364;
  wire seg_2_15_glb_netwk_0_5;
  wire seg_2_15_glb_netwk_4_9;
  wire seg_2_15_local_g0_1_13034;
  wire seg_2_15_local_g0_2_13035;
  wire seg_2_15_local_g0_3_13036;
  wire seg_2_15_local_g0_4_13037;
  wire seg_2_15_local_g0_6_13039;
  wire seg_2_15_local_g0_7_13040;
  wire seg_2_15_local_g1_2_13043;
  wire seg_2_15_local_g2_6_13055;
  wire seg_2_15_local_g3_3_13060;
  wire seg_2_15_local_g3_5_13062;
  wire seg_2_15_local_g3_6_13063;
  wire seg_2_15_lutff_1_out_8773;
  wire seg_2_15_lutff_2_out_8774;
  wire seg_2_15_lutff_3_out_8775;
  wire seg_2_15_lutff_4_out_8776;
  wire seg_2_15_lutff_6_out_8778;
  wire seg_2_15_neigh_op_bnl_6_2819;
  wire seg_2_15_neigh_op_lft_2_3027;
  wire seg_2_15_neigh_op_tnl_3_3253;
  wire seg_2_15_neigh_op_top_1_8920;
  wire seg_2_15_neigh_op_top_2_8921;
  wire seg_2_15_neigh_op_top_6_8925;
  wire seg_2_15_neigh_op_top_7_8926;
  wire seg_2_15_sp4_h_r_10_13129;
  wire seg_2_15_sp4_h_r_14_8936;
  wire seg_2_15_sp4_h_r_29_3341;
  wire seg_2_15_sp4_h_r_30_3342;
  wire seg_2_15_sp4_v_b_19_8656;
  wire seg_2_16_glb_netwk_0_5;
  wire seg_2_16_glb_netwk_4_9;
  wire seg_2_16_local_g0_2_13158;
  wire seg_2_16_local_g0_7_13163;
  wire seg_2_16_local_g1_0_13164;
  wire seg_2_16_local_g1_2_13166;
  wire seg_2_16_local_g2_1_13173;
  wire seg_2_16_local_g2_2_13174;
  wire seg_2_16_local_g3_3_13183;
  wire seg_2_16_local_g3_7_13187;
  wire seg_2_16_lutff_0_out_8919;
  wire seg_2_16_lutff_1_out_8920;
  wire seg_2_16_lutff_2_out_8921;
  wire seg_2_16_lutff_3_out_8922;
  wire seg_2_16_lutff_4_out_8923;
  wire seg_2_16_lutff_5_out_8924;
  wire seg_2_16_lutff_6_out_8925;
  wire seg_2_16_lutff_7_out_8926;
  wire seg_2_16_neigh_op_lft_2_3252;
  wire seg_2_16_neigh_op_rgt_7_13122;
  wire seg_2_16_neigh_op_tnl_1_3457;
  wire seg_2_16_neigh_op_tnl_2_3458;
  wire seg_2_16_neigh_op_top_2_9068;
  wire seg_2_16_neigh_op_top_7_9073;
  wire seg_2_16_sp4_v_b_11_8659;
  wire seg_2_16_sp4_v_b_43_9097;
  wire seg_2_16_sp4_v_b_4_8654;
  wire seg_2_16_sp4_v_b_5_8653;
  wire seg_2_16_sp4_v_b_7_8655;
  wire seg_2_17_glb_netwk_0_5;
  wire seg_2_17_glb_netwk_4_9;
  wire seg_2_17_local_g1_4_13291;
  wire seg_2_17_local_g1_7_13294;
  wire seg_2_17_local_g2_6_13301;
  wire seg_2_17_lutff_2_out_9068;
  wire seg_2_17_lutff_5_out_9071;
  wire seg_2_17_lutff_7_out_9073;
  wire seg_2_17_neigh_op_tnl_6_3670;
  wire seg_2_17_neigh_op_top_4_9217;
  wire seg_2_17_sp4_h_l_39_3731;
  wire seg_2_17_sp4_h_r_7_13382;
  wire seg_2_17_sp4_v_t_39_9387;
  wire seg_2_18_glb_netwk_0_5;
  wire seg_2_18_glb_netwk_4_9;
  wire seg_2_18_local_g0_1_13403;
  wire seg_2_18_local_g0_5_13407;
  wire seg_2_18_local_g0_6_13408;
  wire seg_2_18_local_g0_7_13409;
  wire seg_2_18_local_g2_3_13421;
  wire seg_2_18_lutff_0_out_9213;
  wire seg_2_18_lutff_1_out_9214;
  wire seg_2_18_lutff_4_out_9217;
  wire seg_2_18_lutff_6_out_9219;
  wire seg_2_18_lutff_7_out_9220;
  wire seg_2_18_neigh_op_top_1_9361;
  wire seg_2_18_neigh_op_top_5_9365;
  wire seg_2_18_neigh_op_top_7_9367;
  wire seg_2_18_sp4_h_r_22_9375;
  wire seg_2_18_sp4_r_v_b_35_13395;
  wire seg_2_19_glb_netwk_0_5;
  wire seg_2_19_glb_netwk_4_9;
  wire seg_2_19_local_g0_3_13528;
  wire seg_2_19_local_g0_4_13529;
  wire seg_2_19_local_g0_6_13531;
  wire seg_2_19_local_g1_0_13533;
  wire seg_2_19_local_g1_4_13537;
  wire seg_2_19_local_g1_5_13538;
  wire seg_2_19_local_g1_7_13540;
  wire seg_2_19_lutff_0_out_9360;
  wire seg_2_19_lutff_1_out_9361;
  wire seg_2_19_lutff_4_out_9364;
  wire seg_2_19_lutff_5_out_9365;
  wire seg_2_19_lutff_6_out_9366;
  wire seg_2_19_lutff_7_out_9367;
  wire seg_2_19_neigh_op_lft_0_3873;
  wire seg_2_19_neigh_op_top_3_9510;
  wire seg_2_19_neigh_op_top_4_9511;
  wire seg_2_19_neigh_op_top_5_9512;
  wire seg_2_19_neigh_op_top_7_9514;
  wire seg_2_19_sp4_h_r_12_9520;
  wire seg_2_19_sp4_v_b_6_9097;
  wire seg_2_1_glb_netwk_0_5;
  wire seg_2_1_glb_netwk_4_9;
  wire seg_2_1_local_g0_1_11272;
  wire seg_2_1_local_g0_7_11278;
  wire seg_2_1_local_g1_0_11279;
  wire seg_2_1_local_g1_4_11283;
  wire seg_2_1_local_g2_6_11293;
  wire seg_2_1_local_g2_7_11294;
  wire seg_2_1_local_g3_0_11295;
  wire seg_2_1_local_g3_7_11302;
  wire seg_2_1_lutff_0_out_6673;
  wire seg_2_1_lutff_1_out_6674;
  wire seg_2_1_lutff_3_out_6676;
  wire seg_2_1_lutff_5_out_6678;
  wire seg_2_1_lutff_7_out_6680;
  wire seg_2_1_neigh_op_rgt_6_11235;
  wire seg_2_1_neigh_op_tnl_7_123;
  wire seg_2_1_neigh_op_top_4_6829;
  wire seg_2_1_sp4_r_v_b_0_11381;
  wire seg_2_1_sp4_v_b_42_6886;
  wire seg_2_1_sp4_v_b_47_6891;
  wire seg_2_20_glb_netwk_0_5;
  wire seg_2_20_glb_netwk_4_9;
  wire seg_2_20_local_g0_2_13650;
  wire seg_2_20_local_g0_4_13652;
  wire seg_2_20_local_g0_5_13653;
  wire seg_2_20_local_g0_7_13655;
  wire seg_2_20_local_g3_0_13672;
  wire seg_2_20_lutff_1_out_9508;
  wire seg_2_20_lutff_3_out_9510;
  wire seg_2_20_lutff_4_out_9511;
  wire seg_2_20_lutff_5_out_9512;
  wire seg_2_20_lutff_7_out_9514;
  wire seg_2_20_neigh_op_lft_2_4087;
  wire seg_2_20_neigh_op_tnl_0_4312;
  wire seg_2_20_neigh_op_top_4_9658;
  wire seg_2_20_sp4_h_r_13_9666;
  wire seg_2_20_sp4_v_b_23_9395;
  wire seg_2_20_sp4_v_b_8_9246;
  wire seg_2_21_glb_netwk_0_5;
  wire seg_2_21_glb_netwk_4_9;
  wire seg_2_21_local_g0_5_13776;
  wire seg_2_21_local_g1_0_13779;
  wire seg_2_21_lutff_4_out_9658;
  wire seg_2_21_neigh_op_top_0_9801;
  wire seg_2_21_neigh_op_top_5_9806;
  wire seg_2_21_sp4_v_b_2_9387;
  wire seg_2_21_sp4_v_t_39_9975;
  wire seg_2_22_glb_netwk_0_5;
  wire seg_2_22_glb_netwk_4_9;
  wire seg_2_22_local_g0_3_13897;
  wire seg_2_22_local_g3_2_13920;
  wire seg_2_22_lutff_0_out_9801;
  wire seg_2_22_lutff_5_out_9806;
  wire seg_2_22_neigh_op_tnl_2_4768;
  wire seg_2_22_sp12_h_r_6_4803;
  wire seg_2_22_sp4_h_r_3_13993;
  wire seg_2_22_sp4_v_t_47_10130;
  wire seg_2_23_glb_netwk_0_5;
  wire seg_2_23_glb_netwk_4_9;
  wire seg_2_23_local_g1_1_14026;
  wire seg_2_23_lutff_4_out_9952;
  wire seg_2_23_sp4_h_r_17_10113;
  wire seg_2_24_sp4_v_b_11_9835;
  wire seg_2_25_sp4_h_l_39_5472;
  wire seg_2_25_sp4_h_r_9_14368;
  wire seg_2_26_sp4_h_l_41_5683;
  wire seg_2_2_glb_netwk_0_5;
  wire seg_2_2_glb_netwk_4_9;
  wire seg_2_2_local_g0_1_11435;
  wire seg_2_2_local_g0_2_11436;
  wire seg_2_2_local_g0_3_11437;
  wire seg_2_2_local_g0_4_11438;
  wire seg_2_2_local_g0_5_11439;
  wire seg_2_2_local_g0_6_11440;
  wire seg_2_2_local_g1_0_11442;
  wire seg_2_2_local_g1_2_11444;
  wire seg_2_2_local_g1_3_11445;
  wire seg_2_2_local_g1_4_11446;
  wire seg_2_2_local_g1_5_11447;
  wire seg_2_2_local_g1_6_11448;
  wire seg_2_2_local_g1_7_11449;
  wire seg_2_2_local_g2_1_11451;
  wire seg_2_2_local_g2_2_11452;
  wire seg_2_2_local_g2_4_11454;
  wire seg_2_2_local_g2_5_11455;
  wire seg_2_2_local_g3_4_11462;
  wire seg_2_2_local_g3_7_11465;
  wire seg_2_2_lutff_0_out_6825;
  wire seg_2_2_lutff_1_out_6826;
  wire seg_2_2_lutff_2_out_6827;
  wire seg_2_2_lutff_3_out_6828;
  wire seg_2_2_lutff_4_out_6829;
  wire seg_2_2_lutff_5_out_6830;
  wire seg_2_2_lutff_6_out_6831;
  wire seg_2_2_lutff_7_out_6832;
  wire seg_2_2_neigh_op_bnr_6_11235;
  wire seg_2_2_neigh_op_bot_3_6676;
  wire seg_2_2_neigh_op_bot_5_6678;
  wire seg_2_2_neigh_op_lft_1_117;
  wire seg_2_2_neigh_op_lft_2_118;
  wire seg_2_2_neigh_op_lft_4_120;
  wire seg_2_2_neigh_op_lft_5_121;
  wire seg_2_2_neigh_op_tnl_4_455;
  wire seg_2_2_neigh_op_top_2_7010;
  wire seg_2_2_neigh_op_top_3_7011;
  wire seg_2_2_neigh_op_top_6_7014;
  wire seg_2_2_sp4_h_r_0_11528;
  wire seg_2_2_sp4_h_r_22_7023;
  wire seg_2_2_sp4_h_r_41_523;
  wire seg_2_2_sp4_h_r_47_530;
  wire seg_2_2_sp4_h_r_6_11536;
  wire seg_2_2_sp4_h_r_8_11538;
  wire seg_2_2_sp4_r_v_b_39_11543;
  wire seg_2_2_sp4_v_b_36_7032;
  wire seg_2_2_sp4_v_b_40_7036;
  wire seg_2_2_sp4_v_b_4_6858;
  wire seg_2_2_sp4_v_t_36_7179;
  wire seg_2_3_glb_netwk_0_5;
  wire seg_2_3_glb_netwk_4_9;
  wire seg_2_3_local_g0_1_11558;
  wire seg_2_3_local_g0_3_11560;
  wire seg_2_3_local_g0_4_11561;
  wire seg_2_3_local_g0_5_11562;
  wire seg_2_3_local_g0_6_11563;
  wire seg_2_3_local_g0_7_11564;
  wire seg_2_3_local_g1_0_11565;
  wire seg_2_3_local_g1_2_11567;
  wire seg_2_3_local_g1_4_11569;
  wire seg_2_3_local_g1_5_11570;
  wire seg_2_3_local_g1_7_11572;
  wire seg_2_3_local_g2_0_11573;
  wire seg_2_3_local_g2_2_11575;
  wire seg_2_3_local_g3_4_11585;
  wire seg_2_3_local_g3_5_11586;
  wire seg_2_3_local_g3_7_11588;
  wire seg_2_3_lutff_0_out_7008;
  wire seg_2_3_lutff_1_out_7009;
  wire seg_2_3_lutff_2_out_7010;
  wire seg_2_3_lutff_3_out_7011;
  wire seg_2_3_lutff_4_out_7012;
  wire seg_2_3_lutff_5_out_7013;
  wire seg_2_3_lutff_6_out_7014;
  wire seg_2_3_lutff_7_out_7015;
  wire seg_2_3_neigh_op_bot_0_6825;
  wire seg_2_3_neigh_op_bot_1_6826;
  wire seg_2_3_neigh_op_bot_4_6829;
  wire seg_2_3_neigh_op_bot_6_6831;
  wire seg_2_3_neigh_op_lft_2_453;
  wire seg_2_3_neigh_op_lft_4_455;
  wire seg_2_3_neigh_op_tnr_7_11646;
  wire seg_2_3_neigh_op_top_3_7158;
  wire seg_2_3_neigh_op_top_5_7160;
  wire seg_2_3_sp4_h_l_38_761;
  wire seg_2_3_sp4_h_r_23_7169;
  wire seg_2_3_sp4_r_v_b_21_11421;
  wire seg_2_3_sp4_r_v_b_23_11423;
  wire seg_2_3_sp4_v_b_5_6871;
  wire seg_2_4_glb_netwk_0_5;
  wire seg_2_4_glb_netwk_4_9;
  wire seg_2_4_local_g0_0_11680;
  wire seg_2_4_local_g0_2_11682;
  wire seg_2_4_local_g0_3_11683;
  wire seg_2_4_local_g0_4_11684;
  wire seg_2_4_local_g0_6_11686;
  wire seg_2_4_local_g1_2_11690;
  wire seg_2_4_local_g1_4_11692;
  wire seg_2_4_local_g1_5_11693;
  wire seg_2_4_local_g1_7_11695;
  wire seg_2_4_local_g2_0_11696;
  wire seg_2_4_local_g2_3_11699;
  wire seg_2_4_local_g2_6_11702;
  wire seg_2_4_local_g3_0_11704;
  wire seg_2_4_local_g3_2_11706;
  wire seg_2_4_local_g3_3_11707;
  wire seg_2_4_local_g3_4_11708;
  wire seg_2_4_local_g3_5_11709;
  wire seg_2_4_local_g3_6_11710;
  wire seg_2_4_lutff_0_out_7155;
  wire seg_2_4_lutff_1_out_7156;
  wire seg_2_4_lutff_2_out_7157;
  wire seg_2_4_lutff_3_out_7158;
  wire seg_2_4_lutff_4_out_7159;
  wire seg_2_4_lutff_5_out_7160;
  wire seg_2_4_lutff_6_out_7161;
  wire seg_2_4_lutff_7_out_7162;
  wire seg_2_4_neigh_op_bnl_3_454;
  wire seg_2_4_neigh_op_bnl_5_456;
  wire seg_2_4_neigh_op_bnl_6_457;
  wire seg_2_4_neigh_op_bot_2_7010;
  wire seg_2_4_neigh_op_bot_3_7011;
  wire seg_2_4_neigh_op_lft_2_680;
  wire seg_2_4_neigh_op_lft_4_682;
  wire seg_2_4_neigh_op_lft_5_683;
  wire seg_2_4_neigh_op_lft_7_685;
  wire seg_2_4_neigh_op_rgt_3_11642;
  wire seg_2_4_neigh_op_rgt_4_11643;
  wire seg_2_4_neigh_op_rgt_6_11645;
  wire seg_2_4_neigh_op_tnr_0_11762;
  wire seg_2_4_neigh_op_top_6_7308;
  wire seg_2_4_sp4_h_r_10_11776;
  wire seg_2_4_sp4_v_b_10_6891;
  wire seg_2_4_sp4_v_b_16_7036;
  wire seg_2_4_sp4_v_b_8_6889;
  wire seg_2_5_glb_netwk_0_5;
  wire seg_2_5_glb_netwk_4_9;
  wire seg_2_5_local_g0_6_11809;
  wire seg_2_5_local_g1_5_11816;
  wire seg_2_5_local_g2_0_11819;
  wire seg_2_5_local_g2_2_11821;
  wire seg_2_5_local_g2_6_11825;
  wire seg_2_5_local_g3_2_11829;
  wire seg_2_5_local_g3_4_11831;
  wire seg_2_5_local_g3_6_11833;
  wire seg_2_5_lutff_2_out_7304;
  wire seg_2_5_lutff_4_out_7306;
  wire seg_2_5_lutff_6_out_7308;
  wire seg_2_5_lutff_7_out_7309;
  wire seg_2_5_neigh_op_bnl_2_680;
  wire seg_2_5_neigh_op_lft_6_911;
  wire seg_2_5_neigh_op_rgt_0_11762;
  wire seg_2_5_neigh_op_rgt_4_11766;
  wire seg_2_5_neigh_op_rgt_6_11768;
  wire seg_2_5_sp4_h_l_37_1195;
  wire seg_2_5_sp4_h_l_41_1199;
  wire seg_2_5_sp4_h_l_47_1206;
  wire seg_2_5_sp4_h_r_32_1224;
  wire seg_2_5_sp4_h_r_5_11904;
  wire seg_2_5_sp4_r_v_b_29_11790;
  wire seg_2_5_sp4_r_v_b_39_11912;
  wire seg_2_5_sp4_v_b_12_7179;
  wire seg_2_5_sp4_v_b_32_7335;
  wire seg_2_5_sp4_v_t_39_7623;
  wire seg_2_6_glb_netwk_0_5;
  wire seg_2_6_glb_netwk_4_9;
  wire seg_2_6_local_g0_4_11930;
  wire seg_2_6_local_g1_7_11941;
  wire seg_2_6_local_g2_1_11943;
  wire seg_2_6_local_g3_0_11950;
  wire seg_2_6_local_g3_4_11954;
  wire seg_2_6_local_g3_6_11956;
  wire seg_2_6_local_g3_7_11957;
  wire seg_2_6_lutff_0_out_7449;
  wire seg_2_6_lutff_3_out_7452;
  wire seg_2_6_lutff_4_out_7453;
  wire seg_2_6_lutff_5_out_7454;
  wire seg_2_6_neigh_op_tnr_1_12009;
  wire seg_2_6_neigh_op_tnr_4_12012;
  wire seg_2_6_neigh_op_tnr_6_12014;
  wire seg_2_6_neigh_op_tnr_7_12015;
  wire seg_2_6_sp4_h_r_10_12022;
  wire seg_2_6_sp4_h_r_12_7609;
  wire seg_2_6_sp4_h_r_20_7619;
  wire seg_2_6_sp4_h_r_32_1430;
  wire seg_2_6_sp4_h_r_34_1386;
  wire seg_2_6_sp4_h_r_9_12031;
  wire seg_2_6_sp4_r_v_b_13_11787;
  wire seg_2_6_sp4_r_v_b_21_11795;
  wire seg_2_6_sp4_v_b_15_7329;
  wire seg_2_7_glb_netwk_0_5;
  wire seg_2_7_glb_netwk_3_8;
  wire seg_2_7_local_g0_1_12050;
  wire seg_2_7_local_g0_4_12053;
  wire seg_2_7_local_g0_5_12054;
  wire seg_2_7_local_g0_7_12056;
  wire seg_2_7_local_g2_0_12065;
  wire seg_2_7_local_g2_2_12067;
  wire seg_2_7_local_g2_6_12071;
  wire seg_2_7_local_g3_0_12073;
  wire seg_2_7_local_g3_4_12077;
  wire seg_2_7_lutff_0_out_7596;
  wire seg_2_7_lutff_3_out_7599;
  wire seg_2_7_lutff_4_out_7600;
  wire seg_2_7_lutff_6_out_7602;
  wire seg_2_7_lutff_7_out_7603;
  wire seg_2_7_neigh_op_lft_1_1337;
  wire seg_2_7_sp4_h_l_45_1618;
  wire seg_2_7_sp4_h_r_20_7766;
  wire seg_2_7_sp4_h_r_5_12150;
  wire seg_2_7_sp4_h_r_7_12152;
  wire seg_2_7_sp4_r_v_b_10_11797;
  wire seg_2_7_sp4_r_v_b_3_11788;
  wire seg_2_7_sp4_v_b_30_7627;
  wire seg_2_7_sp4_v_b_36_7767;
  wire seg_2_7_sp4_v_b_40_7771;
  wire seg_2_7_sp4_v_b_8_7335;
  wire seg_2_7_sp4_v_t_37_7915;
  wire seg_2_7_sp4_v_t_42_7920;
  wire seg_2_8_glb_netwk_0_5;
  wire seg_2_8_local_g0_0_12172;
  wire seg_2_8_local_g0_2_12174;
  wire seg_2_8_local_g0_3_12175;
  wire seg_2_8_local_g0_4_12176;
  wire seg_2_8_local_g0_5_12177;
  wire seg_2_8_local_g0_6_12178;
  wire seg_2_8_local_g0_7_12179;
  wire seg_2_8_local_g1_0_12180;
  wire seg_2_8_local_g1_1_12181;
  wire seg_2_8_local_g1_2_12182;
  wire seg_2_8_local_g1_3_12183;
  wire seg_2_8_local_g1_4_12184;
  wire seg_2_8_local_g1_6_12186;
  wire seg_2_8_local_g1_7_12187;
  wire seg_2_8_local_g2_2_12190;
  wire seg_2_8_local_g2_5_12193;
  wire seg_2_8_local_g2_6_12194;
  wire seg_2_8_local_g3_5_12201;
  wire seg_2_8_lutff_2_out_7745;
  wire seg_2_8_lutff_5_out_7748;
  wire seg_2_8_lutff_6_out_7749;
  wire seg_2_8_lutff_7_out_7750;
  wire seg_2_8_neigh_op_bot_3_7599;
  wire seg_2_8_neigh_op_bot_4_7600;
  wire seg_2_8_neigh_op_bot_6_7602;
  wire seg_2_8_neigh_op_bot_7_7603;
  wire seg_2_8_neigh_op_top_6_7896;
  wire seg_2_8_sp4_h_r_0_12266;
  wire seg_2_8_sp4_h_r_18_7911;
  wire seg_2_8_sp4_h_r_1_12267;
  wire seg_2_8_sp4_h_r_2_12270;
  wire seg_2_8_sp4_h_r_3_12271;
  wire seg_2_8_sp4_h_r_6_12274;
  wire seg_2_8_sp4_h_r_8_12276;
  wire seg_2_8_sp4_r_v_b_33_12163;
  wire seg_2_8_sp4_r_v_b_35_12165;
  wire seg_2_8_sp4_v_b_12_7620;
  wire seg_2_8_sp4_v_b_29_7771;
  wire seg_2_8_sp4_v_b_37_7915;
  wire seg_2_8_sp4_v_t_40_8065;
  wire seg_2_9_glb_netwk_0_5;
  wire seg_2_9_glb_netwk_4_9;
  wire seg_2_9_local_g0_0_12295;
  wire seg_2_9_local_g0_2_12297;
  wire seg_2_9_local_g0_4_12299;
  wire seg_2_9_local_g0_5_12300;
  wire seg_2_9_local_g0_7_12302;
  wire seg_2_9_local_g1_5_12308;
  wire seg_2_9_local_g2_1_12312;
  wire seg_2_9_local_g3_0_12319;
  wire seg_2_9_lutff_0_out_7890;
  wire seg_2_9_lutff_1_out_7891;
  wire seg_2_9_lutff_2_out_7892;
  wire seg_2_9_lutff_4_out_7894;
  wire seg_2_9_lutff_5_out_7895;
  wire seg_2_9_lutff_6_out_7896;
  wire seg_2_9_neigh_op_lft_5_1758;
  wire seg_2_9_neigh_op_lft_7_1760;
  wire seg_2_9_neigh_op_tnl_1_1966;
  wire seg_2_9_sp12_h_r_12_2012;
  wire seg_2_9_sp4_h_r_0_12389;
  wire seg_2_9_sp4_h_r_12_8050;
  wire seg_2_9_sp4_h_r_22_8052;
  wire seg_2_9_sp4_h_r_8_12399;
  wire seg_2_9_sp4_r_v_b_13_12156;
  wire seg_2_9_sp4_r_v_b_23_12166;
  wire seg_2_9_sp4_r_v_b_31_12284;
  wire seg_2_9_sp4_r_v_b_39_12404;
  wire seg_2_9_sp4_v_b_12_7767;
  wire seg_2_9_sp4_v_b_21_7776;
  wire seg_2_9_sp4_v_b_32_7923;
  wire seg_2_9_sp4_v_b_3_7622;
  wire seg_2_9_sp4_v_b_46_8071;
  wire seg_2_9_sp4_v_b_4_7625;
  wire seg_2_9_sp4_v_b_5_7624;
  wire seg_2_9_sp4_v_t_43_8215;
  wire seg_2_9_sp4_v_t_47_8219;
  wire seg_3_10_glb_netwk_0_5;
  wire seg_3_10_glb_netwk_4_9;
  wire seg_3_10_local_g0_4_16253;
  wire seg_3_10_local_g0_5_16254;
  wire seg_3_10_local_g1_3_16260;
  wire seg_3_10_local_g1_4_16261;
  wire seg_3_10_local_g2_3_16268;
  wire seg_3_10_local_g3_0_16273;
  wire seg_3_10_local_g3_3_16276;
  wire seg_3_10_local_g3_5_16278;
  wire seg_3_10_lutff_0_out_12377;
  wire seg_3_10_lutff_1_out_12378;
  wire seg_3_10_lutff_3_out_12380;
  wire seg_3_10_lutff_4_out_12381;
  wire seg_3_10_lutff_5_out_12382;
  wire seg_3_10_lutff_7_out_12384;
  wire seg_3_10_neigh_op_top_4_12504;
  wire seg_3_10_sp4_h_l_42_2248;
  wire seg_3_10_sp4_h_r_11_16346;
  wire seg_3_10_sp4_h_r_13_12512;
  wire seg_3_10_sp4_h_r_19_12520;
  wire seg_3_10_sp4_h_r_20_12523;
  wire seg_3_10_sp4_h_r_43_2282;
  wire seg_3_10_sp4_h_r_4_16349;
  wire seg_3_10_sp4_h_r_7_16352;
  wire seg_3_10_sp4_h_r_9_16354;
  wire seg_3_10_sp4_r_v_b_29_16236;
  wire seg_3_10_sp4_v_b_0_12156;
  wire seg_3_10_sp4_v_b_10_12166;
  wire seg_3_10_sp4_v_b_11_12165;
  wire seg_3_10_sp4_v_b_27_12403;
  wire seg_3_10_sp4_v_b_32_12410;
  wire seg_3_10_sp4_v_b_4_12160;
  wire seg_3_10_sp4_v_b_8_12164;
  wire seg_3_10_sp4_v_b_9_12163;
  wire seg_3_10_sp4_v_t_43_12654;
  wire seg_3_11_glb_netwk_0_5;
  wire seg_3_11_glb_netwk_4_9;
  wire seg_3_11_local_g0_3_16375;
  wire seg_3_11_local_g1_3_16383;
  wire seg_3_11_local_g1_5_16385;
  wire seg_3_11_local_g1_6_16386;
  wire seg_3_11_local_g1_7_16387;
  wire seg_3_11_local_g2_0_16388;
  wire seg_3_11_local_g2_2_16390;
  wire seg_3_11_local_g2_6_16394;
  wire seg_3_11_lutff_2_out_12502;
  wire seg_3_11_lutff_4_out_12504;
  wire seg_3_11_lutff_7_out_12507;
  wire seg_3_11_neigh_op_lft_5_8189;
  wire seg_3_11_sp4_h_l_36_2448;
  wire seg_3_11_sp4_h_r_11_16469;
  wire seg_3_11_sp4_h_r_14_12640;
  wire seg_3_11_sp4_h_r_15_12639;
  wire seg_3_11_sp4_h_r_3_16471;
  wire seg_3_11_sp4_h_r_42_2489;
  wire seg_3_11_sp4_h_r_44_2491;
  wire seg_3_11_sp4_h_r_8_16476;
  wire seg_3_11_sp4_r_v_b_14_16234;
  wire seg_3_11_sp4_r_v_b_1_16109;
  wire seg_3_11_sp4_r_v_b_27_16357;
  wire seg_3_11_sp4_r_v_b_29_16359;
  wire seg_3_11_sp4_r_v_b_33_16363;
  wire seg_3_11_sp4_r_v_b_3_16111;
  wire seg_3_11_sp4_r_v_b_7_16115;
  wire seg_3_11_sp4_v_b_11_12288;
  wire seg_3_11_sp4_v_b_18_12407;
  wire seg_3_11_sp4_v_b_22_12411;
  wire seg_3_11_sp4_v_b_32_12533;
  wire seg_3_11_sp4_v_b_6_12285;
  wire seg_3_11_sp4_v_b_7_12284;
  wire seg_3_12_local_g0_3_16498;
  wire seg_3_12_local_g0_4_16499;
  wire seg_3_12_local_g0_5_16500;
  wire seg_3_12_local_g1_1_16504;
  wire seg_3_12_local_g1_4_16507;
  wire seg_3_12_local_g1_5_16508;
  wire seg_3_12_local_g1_7_16510;
  wire seg_3_12_local_g2_2_16513;
  wire seg_3_12_local_g2_3_16514;
  wire seg_3_12_local_g2_4_16515;
  wire seg_3_12_local_g2_6_16517;
  wire seg_3_12_local_g2_7_16518;
  wire seg_3_12_local_g3_4_16523;
  wire seg_3_12_local_g3_6_16525;
  wire seg_3_12_lutff_1_out_12624;
  wire seg_3_12_lutff_2_out_12625;
  wire seg_3_12_lutff_3_out_12626;
  wire seg_3_12_lutff_4_out_12627;
  wire seg_3_12_lutff_5_out_12628;
  wire seg_3_12_lutff_6_out_12629;
  wire seg_3_12_lutff_7_out_12630;
  wire seg_3_12_neigh_op_bot_7_12507;
  wire seg_3_12_neigh_op_rgt_2_16456;
  wire seg_3_12_neigh_op_tnl_4_8482;
  wire seg_3_12_neigh_op_tnl_6_8484;
  wire seg_3_12_sp4_h_l_37_2657;
  wire seg_3_12_sp4_h_l_40_2660;
  wire seg_3_12_sp4_h_l_44_2665;
  wire seg_3_12_sp4_h_r_10_16591;
  wire seg_3_12_sp4_h_r_12_12759;
  wire seg_3_12_sp4_h_r_13_12758;
  wire seg_3_12_sp4_h_r_1_16590;
  wire seg_3_12_sp4_h_r_3_16594;
  wire seg_3_12_sp4_h_r_4_16595;
  wire seg_3_12_sp4_r_v_b_39_16604;
  wire seg_3_12_sp4_v_b_0_12402;
  wire seg_3_12_sp4_v_b_11_12411;
  wire seg_3_12_sp4_v_b_13_12525;
  wire seg_3_12_sp4_v_b_2_12404;
  wire seg_3_12_sp4_v_b_35_12657;
  wire seg_3_12_sp4_v_b_36_12770;
  wire seg_3_12_sp4_v_b_46_12780;
  wire seg_3_12_sp4_v_b_7_12407;
  wire seg_3_12_sp4_v_t_37_12894;
  wire seg_3_12_sp4_v_t_42_12899;
  wire seg_3_12_sp4_v_t_43_12900;
  wire seg_3_12_sp4_v_t_46_12903;
  wire seg_3_13_glb_netwk_0_5;
  wire seg_3_13_glb_netwk_4_9;
  wire seg_3_13_local_g0_5_16623;
  wire seg_3_13_local_g0_7_16625;
  wire seg_3_13_local_g1_7_16633;
  wire seg_3_13_local_g2_0_16634;
  wire seg_3_13_local_g2_2_16636;
  wire seg_3_13_local_g2_3_16637;
  wire seg_3_13_local_g2_4_16638;
  wire seg_3_13_local_g2_5_16639;
  wire seg_3_13_local_g2_6_16640;
  wire seg_3_13_local_g3_0_16642;
  wire seg_3_13_local_g3_1_16643;
  wire seg_3_13_local_g3_2_16644;
  wire seg_3_13_local_g3_3_16645;
  wire seg_3_13_local_g3_4_16646;
  wire seg_3_13_local_g3_5_16647;
  wire seg_3_13_local_g3_6_16648;
  wire seg_3_13_lutff_7_out_12753;
  wire seg_3_13_neigh_op_bnl_0_8331;
  wire seg_3_13_neigh_op_bnl_1_8332;
  wire seg_3_13_neigh_op_bnl_2_8333;
  wire seg_3_13_neigh_op_bnl_3_8334;
  wire seg_3_13_neigh_op_bnl_4_8335;
  wire seg_3_13_neigh_op_bnl_5_8336;
  wire seg_3_13_neigh_op_bnl_6_8337;
  wire seg_3_13_neigh_op_top_5_12874;
  wire seg_3_13_sp4_h_l_39_2868;
  wire seg_3_13_sp4_h_l_41_2870;
  wire seg_3_13_sp4_h_l_43_2872;
  wire seg_3_13_sp4_h_r_10_16714;
  wire seg_3_13_sp4_h_r_12_12882;
  wire seg_3_13_sp4_h_r_20_12892;
  wire seg_3_13_sp4_h_r_22_12884;
  wire seg_3_13_sp4_h_r_2_16716;
  wire seg_3_13_sp4_h_r_7_16721;
  wire seg_3_13_sp4_h_r_8_16722;
  wire seg_3_13_sp4_r_v_b_31_16607;
  wire seg_3_13_sp4_r_v_b_37_16725;
  wire seg_3_13_sp4_r_v_b_43_16731;
  wire seg_3_13_sp4_v_b_28_12775;
  wire seg_3_13_sp4_v_b_32_12779;
  wire seg_3_13_sp4_v_b_34_12781;
  wire seg_3_13_sp4_v_b_38_12895;
  wire seg_3_13_sp4_v_b_7_12530;
  wire seg_3_13_sp4_v_t_36_13016;
  wire seg_3_13_sp4_v_t_37_13017;
  wire seg_3_13_sp4_v_t_38_13018;
  wire seg_3_14_glb_netwk_0_5;
  wire seg_3_14_glb_netwk_4_9;
  wire seg_3_14_local_g0_1_16742;
  wire seg_3_14_local_g0_7_16748;
  wire seg_3_14_local_g1_7_16756;
  wire seg_3_14_local_g2_0_16757;
  wire seg_3_14_local_g2_1_16758;
  wire seg_3_14_local_g2_4_16761;
  wire seg_3_14_local_g2_5_16762;
  wire seg_3_14_local_g3_0_16765;
  wire seg_3_14_local_g3_2_16767;
  wire seg_3_14_local_g3_3_16768;
  wire seg_3_14_local_g3_5_16770;
  wire seg_3_14_lutff_0_out_12869;
  wire seg_3_14_lutff_1_out_12870;
  wire seg_3_14_lutff_2_out_12871;
  wire seg_3_14_lutff_5_out_12874;
  wire seg_3_14_neigh_op_bnl_0_8478;
  wire seg_3_14_neigh_op_rgt_0_16700;
  wire seg_3_14_neigh_op_rgt_3_16703;
  wire seg_3_14_neigh_op_tnr_5_16828;
  wire seg_3_14_neigh_op_top_7_12999;
  wire seg_3_14_sp4_h_l_36_3092;
  wire seg_3_14_sp4_r_v_b_15_16604;
  wire seg_3_14_sp4_v_b_0_12648;
  wire seg_3_14_sp4_v_b_12_12770;
  wire seg_3_14_sp4_v_b_1_12647;
  wire seg_3_14_sp4_v_b_24_12894;
  wire seg_3_14_sp4_v_b_25_12893;
  wire seg_3_14_sp4_v_b_28_12898;
  wire seg_3_14_sp4_v_b_29_12897;
  wire seg_3_14_sp4_v_b_2_12650;
  wire seg_3_14_sp4_v_b_6_12654;
  wire seg_3_14_sp4_v_b_7_12653;
  wire seg_3_14_sp4_v_b_8_12656;
  wire seg_3_14_sp4_v_b_9_12655;
  wire seg_3_14_sp4_v_t_45_13148;
  wire seg_3_15_local_g0_0_16864;
  wire seg_3_15_local_g0_2_16866;
  wire seg_3_15_local_g0_3_16867;
  wire seg_3_15_local_g0_4_16868;
  wire seg_3_15_local_g0_5_16869;
  wire seg_3_15_local_g1_1_16873;
  wire seg_3_15_local_g1_6_16878;
  wire seg_3_15_local_g2_3_16883;
  wire seg_3_15_local_g2_4_16884;
  wire seg_3_15_local_g2_6_16886;
  wire seg_3_15_local_g3_2_16890;
  wire seg_3_15_local_g3_4_16892;
  wire seg_3_15_local_g3_5_16893;
  wire seg_3_15_local_g3_6_16894;
  wire seg_3_15_lutff_7_out_12999;
  wire seg_3_15_neigh_op_bnr_3_16703;
  wire seg_3_15_neigh_op_lft_6_8778;
  wire seg_3_15_neigh_op_rgt_2_16825;
  wire seg_3_15_neigh_op_rgt_3_16826;
  wire seg_3_15_neigh_op_rgt_4_16827;
  wire seg_3_15_neigh_op_tnl_4_8923;
  wire seg_3_15_neigh_op_tnl_5_8924;
  wire seg_3_15_neigh_op_tnr_6_16952;
  wire seg_3_15_neigh_op_top_0_13115;
  wire seg_3_15_neigh_op_top_1_13116;
  wire seg_3_15_neigh_op_top_2_13117;
  wire seg_3_15_neigh_op_top_4_13119;
  wire seg_3_15_neigh_op_top_5_13120;
  wire seg_3_15_sp4_h_l_38_3304;
  wire seg_3_15_sp4_h_l_40_3306;
  wire seg_3_15_sp4_h_l_42_3308;
  wire seg_3_15_sp4_h_r_4_16964;
  wire seg_3_15_sp4_r_v_b_13_16725;
  wire seg_3_15_sp4_r_v_b_19_16731;
  wire seg_3_15_sp4_r_v_b_7_16607;
  wire seg_3_15_sp4_v_b_10_12781;
  wire seg_3_15_sp4_v_b_14_12895;
  wire seg_3_15_sp4_v_b_38_13141;
  wire seg_3_15_sp4_v_b_4_12775;
  wire seg_3_15_sp4_v_b_7_12776;
  wire seg_3_15_sp4_v_b_8_12779;
  wire seg_3_15_sp4_v_b_9_12778;
  wire seg_3_15_sp4_v_t_38_13264;
  wire seg_3_16_glb_netwk_0_5;
  wire seg_3_16_glb_netwk_4_9;
  wire seg_3_16_local_g0_2_16989;
  wire seg_3_16_local_g0_3_16990;
  wire seg_3_16_local_g0_5_16992;
  wire seg_3_16_local_g1_3_16998;
  wire seg_3_16_local_g1_4_16999;
  wire seg_3_16_local_g1_6_17001;
  wire seg_3_16_local_g2_1_17004;
  wire seg_3_16_local_g3_5_17016;
  wire seg_3_16_lutff_0_out_13115;
  wire seg_3_16_lutff_1_out_13116;
  wire seg_3_16_lutff_2_out_13117;
  wire seg_3_16_lutff_4_out_13119;
  wire seg_3_16_lutff_5_out_13120;
  wire seg_3_16_lutff_7_out_13122;
  wire seg_3_16_neigh_op_lft_3_8922;
  wire seg_3_16_neigh_op_rgt_1_16947;
  wire seg_3_16_neigh_op_tnl_5_9071;
  wire seg_3_16_neigh_op_top_2_13240;
  wire seg_3_16_neigh_op_top_3_13241;
  wire seg_3_16_neigh_op_top_4_13242;
  wire seg_3_16_neigh_op_top_5_13243;
  wire seg_3_16_neigh_op_top_6_13244;
  wire seg_3_16_sp4_h_l_42_3514;
  wire seg_3_16_sp4_v_b_10_12904;
  wire seg_3_16_sp4_v_b_12_13016;
  wire seg_3_16_sp4_v_b_2_12896;
  wire seg_3_16_sp4_v_b_4_12898;
  wire seg_3_16_sp4_v_b_6_12900;
  wire seg_3_16_sp4_v_t_39_13388;
  wire seg_3_17_glb_netwk_0_5;
  wire seg_3_17_glb_netwk_4_9;
  wire seg_3_17_local_g0_4_17114;
  wire seg_3_17_local_g0_5_17115;
  wire seg_3_17_local_g1_3_17121;
  wire seg_3_17_local_g2_0_17126;
  wire seg_3_17_local_g2_1_17127;
  wire seg_3_17_local_g2_6_17132;
  wire seg_3_17_local_g2_7_17133;
  wire seg_3_17_lutff_2_out_13240;
  wire seg_3_17_lutff_3_out_13241;
  wire seg_3_17_lutff_4_out_13242;
  wire seg_3_17_lutff_5_out_13243;
  wire seg_3_17_lutff_6_out_13244;
  wire seg_3_17_neigh_op_tnl_0_9213;
  wire seg_3_17_neigh_op_tnl_1_9214;
  wire seg_3_17_neigh_op_tnl_6_9219;
  wire seg_3_17_neigh_op_tnl_7_9220;
  wire seg_3_17_sp4_h_r_10_17206;
  wire seg_3_17_sp4_h_r_3_17209;
  wire seg_3_17_sp4_r_v_b_29_17097;
  wire seg_3_17_sp4_v_b_0_13017;
  wire seg_3_17_sp4_v_b_12_13139;
  wire seg_3_17_sp4_v_b_14_13141;
  wire seg_3_17_sp4_v_b_7_13022;
  wire seg_3_17_sp4_v_t_47_13519;
  wire seg_3_18_glb_netwk_0_5;
  wire seg_3_18_glb_netwk_4_9;
  wire seg_3_18_local_g0_0_17233;
  wire seg_3_18_local_g0_1_17234;
  wire seg_3_18_local_g0_4_17237;
  wire seg_3_18_local_g0_5_17238;
  wire seg_3_18_local_g1_0_17241;
  wire seg_3_18_local_g1_1_17242;
  wire seg_3_18_local_g1_2_17243;
  wire seg_3_18_local_g1_3_17244;
  wire seg_3_18_local_g1_4_17245;
  wire seg_3_18_local_g1_5_17246;
  wire seg_3_18_local_g1_7_17248;
  wire seg_3_18_local_g2_0_17249;
  wire seg_3_18_local_g2_4_17253;
  wire seg_3_18_local_g3_2_17259;
  wire seg_3_18_neigh_op_tnl_4_9364;
  wire seg_3_18_neigh_op_top_5_13489;
  wire seg_3_18_sp4_r_v_b_11_16980;
  wire seg_3_18_sp4_r_v_b_13_17094;
  wire seg_3_18_sp4_r_v_b_18_17099;
  wire seg_3_18_sp4_r_v_b_1_16970;
  wire seg_3_18_sp4_r_v_b_2_16973;
  wire seg_3_18_sp4_r_v_b_3_16972;
  wire seg_3_18_sp4_r_v_b_4_16975;
  wire seg_3_18_sp4_r_v_b_8_16979;
  wire seg_3_18_sp4_v_b_0_13140;
  wire seg_3_18_sp4_v_b_14_13264;
  wire seg_3_18_sp4_v_b_16_13266;
  wire seg_3_18_sp4_v_b_17_13267;
  wire seg_3_18_sp4_v_b_23_13273;
  wire seg_3_18_sp4_v_b_4_13144;
  wire seg_3_18_sp4_v_b_5_13143;
  wire seg_3_18_sp4_v_b_8_13148;
  wire seg_3_18_sp4_v_b_9_13147;
  wire seg_3_18_sp4_v_t_36_13631;
  wire seg_3_19_glb_netwk_0_5;
  wire seg_3_19_glb_netwk_4_9;
  wire seg_3_19_local_g1_0_17364;
  wire seg_3_19_local_g2_1_17373;
  wire seg_3_19_lutff_5_out_13489;
  wire seg_3_19_neigh_op_lft_0_9360;
  wire seg_3_19_neigh_op_tnl_1_9508;
  wire seg_3_19_sp4_r_v_b_5_17097;
  wire seg_3_1_glb_netwk_0_5;
  wire seg_3_1_glb_netwk_4_9;
  wire seg_3_1_local_g0_1_15103;
  wire seg_3_1_local_g0_2_15104;
  wire seg_3_1_local_g0_4_15106;
  wire seg_3_1_local_g1_0_15110;
  wire seg_3_1_local_g1_5_15115;
  wire seg_3_1_local_g2_0_15118;
  wire seg_3_1_local_g2_1_15119;
  wire seg_3_1_local_g2_2_15120;
  wire seg_3_1_local_g2_3_15121;
  wire seg_3_1_local_g2_4_15122;
  wire seg_3_1_local_g2_6_15124;
  wire seg_3_1_local_g3_0_15126;
  wire seg_3_1_local_g3_1_15127;
  wire seg_3_1_local_g3_3_15129;
  wire seg_3_1_local_g3_5_15131;
  wire seg_3_1_local_g3_6_15132;
  wire seg_3_1_local_g3_7_15133;
  wire seg_3_1_lutff_0_out_11229;
  wire seg_3_1_lutff_1_out_11230;
  wire seg_3_1_lutff_2_out_11231;
  wire seg_3_1_lutff_3_out_11232;
  wire seg_3_1_lutff_6_out_11235;
  wire seg_3_1_lutff_7_out_11236;
  wire seg_3_1_neigh_op_rgt_0_15060;
  wire seg_3_1_neigh_op_rgt_3_15063;
  wire seg_3_1_neigh_op_rgt_5_15065;
  wire seg_3_1_neigh_op_rgt_6_15066;
  wire seg_3_1_neigh_op_rgt_7_15067;
  wire seg_3_1_neigh_op_tnl_3_6828;
  wire seg_3_1_neigh_op_tnr_6_15194;
  wire seg_3_1_sp4_h_r_12_11370;
  wire seg_3_1_sp4_h_r_13_11369;
  wire seg_3_1_sp4_h_r_14_11374;
  wire seg_3_1_sp4_h_r_16_11376;
  wire seg_3_1_sp4_h_r_18_11378;
  wire seg_3_1_sp4_h_r_20_11380;
  wire seg_3_1_sp4_h_r_28_6843;
  wire seg_3_1_sp4_h_r_2_15204;
  wire seg_3_1_sp4_h_r_34_6839;
  wire seg_3_1_sp4_h_r_44_250;
  wire seg_3_1_sp4_h_r_4_15206;
  wire seg_3_1_sp4_h_r_6_15208;
  wire seg_3_1_sp4_r_v_b_29_15234;
  wire seg_3_1_sp4_v_b_41_11417;
  wire seg_3_1_sp4_v_t_37_11541;
  wire seg_3_1_sp4_v_t_44_11548;
  wire seg_3_20_glb_netwk_0_5;
  wire seg_3_20_glb_netwk_4_9;
  wire seg_3_20_local_g3_1_17504;
  wire seg_3_20_sp4_h_r_33_9677;
  wire seg_3_20_sp4_v_b_2_13388;
  wire seg_3_20_sp4_v_b_5_13389;
  wire seg_3_20_sp4_v_b_6_13392;
  wire seg_3_20_sp4_v_t_46_13887;
  wire seg_3_21_glb_netwk_0_5;
  wire seg_3_21_glb_netwk_4_9;
  wire seg_3_21_local_g1_3_17613;
  wire seg_3_21_local_g2_2_17620;
  wire seg_3_21_neigh_op_top_3_13856;
  wire seg_3_21_sp4_h_r_26_9817;
  wire seg_3_21_sp4_v_b_10_13519;
  wire seg_3_21_sp4_v_b_12_13631;
  wire seg_3_22_glb_netwk_0_5;
  wire seg_3_22_glb_netwk_4_9;
  wire seg_3_22_local_g2_4_17745;
  wire seg_3_22_lutff_3_out_13856;
  wire seg_3_22_neigh_op_tnl_4_9952;
  wire seg_3_24_sp4_h_l_46_5260;
  wire seg_3_24_sp4_v_b_2_13880;
  wire seg_3_24_sp4_v_b_8_13886;
  wire seg_3_2_glb_netwk_0_5;
  wire seg_3_2_glb_netwk_4_9;
  wire seg_3_2_local_g0_0_15265;
  wire seg_3_2_local_g0_3_15268;
  wire seg_3_2_local_g0_4_15269;
  wire seg_3_2_local_g0_5_15270;
  wire seg_3_2_local_g1_0_15273;
  wire seg_3_2_local_g1_1_15274;
  wire seg_3_2_local_g1_6_15279;
  wire seg_3_2_local_g1_7_15280;
  wire seg_3_2_local_g2_1_15282;
  wire seg_3_2_local_g2_2_15283;
  wire seg_3_2_local_g2_3_15284;
  wire seg_3_2_local_g2_4_15285;
  wire seg_3_2_local_g2_5_15286;
  wire seg_3_2_local_g3_0_15289;
  wire seg_3_2_local_g3_1_15290;
  wire seg_3_2_local_g3_2_15291;
  wire seg_3_2_local_g3_3_15292;
  wire seg_3_2_local_g3_4_15293;
  wire seg_3_2_local_g3_5_15294;
  wire seg_3_2_local_g3_6_15295;
  wire seg_3_2_local_g3_7_15296;
  wire seg_3_2_lutff_0_out_11357;
  wire seg_3_2_lutff_1_out_11358;
  wire seg_3_2_lutff_2_out_11359;
  wire seg_3_2_lutff_3_out_11360;
  wire seg_3_2_lutff_4_out_11361;
  wire seg_3_2_lutff_5_out_11362;
  wire seg_3_2_lutff_6_out_11363;
  wire seg_3_2_lutff_7_out_11364;
  wire seg_3_2_neigh_op_bnr_3_15063;
  wire seg_3_2_neigh_op_rgt_1_15189;
  wire seg_3_2_neigh_op_rgt_4_15192;
  wire seg_3_2_neigh_op_rgt_5_15193;
  wire seg_3_2_neigh_op_top_0_11516;
  wire seg_3_2_sp4_h_r_25_7021;
  wire seg_3_2_sp4_h_r_4_15365;
  wire seg_3_2_sp4_h_r_7_15368;
  wire seg_3_2_sp4_h_r_8_15369;
  wire seg_3_2_sp4_r_v_b_13_15229;
  wire seg_3_2_sp4_r_v_b_24_15243;
  wire seg_3_2_sp4_r_v_b_29_15247;
  wire seg_3_2_sp4_r_v_b_31_15249;
  wire seg_3_2_sp4_r_v_b_34_15254;
  wire seg_3_2_sp4_r_v_b_43_15378;
  wire seg_3_2_sp4_r_v_b_44_15379;
  wire seg_3_2_sp4_v_b_22_11410;
  wire seg_3_2_sp4_v_t_41_11668;
  wire seg_3_3_glb_netwk_0_5;
  wire seg_3_3_glb_netwk_4_9;
  wire seg_3_3_local_g0_2_15390;
  wire seg_3_3_local_g0_3_15391;
  wire seg_3_3_local_g0_4_15392;
  wire seg_3_3_local_g0_6_15394;
  wire seg_3_3_local_g0_7_15395;
  wire seg_3_3_local_g1_1_15397;
  wire seg_3_3_local_g1_2_15398;
  wire seg_3_3_local_g1_3_15399;
  wire seg_3_3_local_g1_4_15400;
  wire seg_3_3_local_g1_6_15402;
  wire seg_3_3_local_g2_0_15404;
  wire seg_3_3_local_g2_2_15406;
  wire seg_3_3_local_g2_3_15407;
  wire seg_3_3_local_g2_4_15408;
  wire seg_3_3_local_g2_5_15409;
  wire seg_3_3_local_g2_6_15410;
  wire seg_3_3_local_g3_0_15412;
  wire seg_3_3_local_g3_2_15414;
  wire seg_3_3_local_g3_3_15415;
  wire seg_3_3_local_g3_4_15416;
  wire seg_3_3_local_g3_5_15417;
  wire seg_3_3_lutff_0_out_11516;
  wire seg_3_3_lutff_1_out_11517;
  wire seg_3_3_lutff_2_out_11518;
  wire seg_3_3_lutff_3_out_11519;
  wire seg_3_3_lutff_4_out_11520;
  wire seg_3_3_lutff_5_out_11521;
  wire seg_3_3_lutff_6_out_11522;
  wire seg_3_3_lutff_7_out_11523;
  wire seg_3_3_neigh_op_bot_6_11363;
  wire seg_3_3_neigh_op_rgt_0_15347;
  wire seg_3_3_neigh_op_rgt_2_15349;
  wire seg_3_3_neigh_op_rgt_3_15350;
  wire seg_3_3_neigh_op_rgt_4_15351;
  wire seg_3_3_neigh_op_tnr_0_15470;
  wire seg_3_3_neigh_op_tnr_3_15473;
  wire seg_3_3_neigh_op_top_2_11641;
  wire seg_3_3_sp4_h_r_11_15485;
  wire seg_3_3_sp4_h_r_20_11662;
  wire seg_3_3_sp4_h_r_26_7171;
  wire seg_3_3_sp4_h_r_29_7174;
  wire seg_3_3_sp4_h_r_4_15488;
  wire seg_3_3_sp4_h_r_6_15490;
  wire seg_3_3_sp4_r_v_b_14_15244;
  wire seg_3_3_sp4_r_v_b_28_15376;
  wire seg_3_3_sp4_v_b_40_11667;
  wire seg_3_3_sp4_v_t_40_11790;
  wire seg_3_4_glb_netwk_0_5;
  wire seg_3_4_glb_netwk_4_9;
  wire seg_3_4_local_g0_0_15511;
  wire seg_3_4_local_g0_3_15514;
  wire seg_3_4_local_g0_5_15516;
  wire seg_3_4_local_g0_7_15518;
  wire seg_3_4_local_g1_0_15519;
  wire seg_3_4_local_g1_3_15522;
  wire seg_3_4_local_g1_4_15523;
  wire seg_3_4_local_g1_5_15524;
  wire seg_3_4_local_g1_6_15525;
  wire seg_3_4_local_g1_7_15526;
  wire seg_3_4_local_g2_0_15527;
  wire seg_3_4_local_g2_3_15530;
  wire seg_3_4_local_g2_6_15533;
  wire seg_3_4_local_g3_1_15536;
  wire seg_3_4_lutff_0_out_11639;
  wire seg_3_4_lutff_2_out_11641;
  wire seg_3_4_lutff_3_out_11642;
  wire seg_3_4_lutff_4_out_11643;
  wire seg_3_4_lutff_5_out_11644;
  wire seg_3_4_lutff_6_out_11645;
  wire seg_3_4_lutff_7_out_11646;
  wire seg_3_4_neigh_op_bnl_1_7009;
  wire seg_3_4_neigh_op_lft_5_7160;
  wire seg_3_4_neigh_op_lft_6_7161;
  wire seg_3_4_neigh_op_lft_7_7162;
  wire seg_3_4_neigh_op_rgt_0_15470;
  wire seg_3_4_neigh_op_rgt_3_15473;
  wire seg_3_4_neigh_op_top_0_11762;
  wire seg_3_4_sp4_h_r_11_15608;
  wire seg_3_4_sp4_h_r_12_11775;
  wire seg_3_4_sp4_h_r_1_15606;
  wire seg_3_4_sp4_h_r_30_7322;
  wire seg_3_4_sp4_h_r_6_15613;
  wire seg_3_4_sp4_r_v_b_1_15242;
  wire seg_3_4_sp4_r_v_b_5_15247;
  wire seg_3_4_sp4_v_b_10_11423;
  wire seg_3_4_sp4_v_b_15_11543;
  wire seg_3_4_sp4_v_b_19_11547;
  wire seg_3_4_sp4_v_b_20_11548;
  wire seg_3_4_sp4_v_b_28_11668;
  wire seg_3_4_sp4_v_b_32_11672;
  wire seg_3_4_sp4_v_b_4_11417;
  wire seg_3_4_sp4_v_b_8_11421;
  wire seg_3_4_sp4_v_t_39_11912;
  wire seg_3_5_glb_netwk_0_5;
  wire seg_3_5_glb_netwk_4_9;
  wire seg_3_5_local_g0_4_15638;
  wire seg_3_5_local_g0_6_15640;
  wire seg_3_5_local_g1_0_15642;
  wire seg_3_5_local_g1_2_15644;
  wire seg_3_5_local_g1_6_15648;
  wire seg_3_5_local_g2_1_15651;
  wire seg_3_5_local_g2_3_15653;
  wire seg_3_5_local_g2_5_15655;
  wire seg_3_5_local_g3_2_15660;
  wire seg_3_5_lutff_0_out_11762;
  wire seg_3_5_lutff_2_out_11764;
  wire seg_3_5_lutff_4_out_11766;
  wire seg_3_5_lutff_6_out_11768;
  wire seg_3_5_neigh_op_bot_0_11639;
  wire seg_3_5_neigh_op_rgt_3_15596;
  wire seg_3_5_neigh_op_tnl_5_7454;
  wire seg_3_5_sp4_h_l_38_1184;
  wire seg_3_5_sp4_h_r_10_15730;
  wire seg_3_5_sp4_h_r_12_11898;
  wire seg_3_5_sp4_h_r_14_11902;
  wire seg_3_5_sp4_h_r_26_7465;
  wire seg_3_5_sp4_h_r_30_7469;
  wire seg_3_5_sp4_h_r_32_7471;
  wire seg_3_5_sp4_h_r_34_7463;
  wire seg_3_5_sp4_h_r_6_15736;
  wire seg_3_5_sp4_r_v_b_18_15500;
  wire seg_3_5_sp4_r_v_b_33_15625;
  wire seg_3_5_sp4_v_b_0_11541;
  wire seg_3_5_sp4_v_b_33_11794;
  wire seg_3_5_sp4_v_t_43_12039;
  wire seg_3_6_glb_netwk_0_5;
  wire seg_3_6_local_g0_4_15761;
  wire seg_3_6_local_g0_5_15762;
  wire seg_3_6_local_g1_0_15765;
  wire seg_3_6_local_g1_1_15766;
  wire seg_3_6_local_g1_2_15767;
  wire seg_3_6_local_g1_5_15770;
  wire seg_3_6_local_g1_7_15772;
  wire seg_3_6_local_g2_1_15774;
  wire seg_3_6_local_g2_2_15775;
  wire seg_3_6_local_g2_3_15776;
  wire seg_3_6_local_g3_0_15781;
  wire seg_3_6_local_g3_2_15783;
  wire seg_3_6_local_g3_3_15784;
  wire seg_3_6_lutff_0_out_11885;
  wire seg_3_6_lutff_1_out_11886;
  wire seg_3_6_lutff_5_out_11890;
  wire seg_3_6_lutff_7_out_11892;
  wire seg_3_6_neigh_op_bnr_5_15598;
  wire seg_3_6_neigh_op_rgt_0_15716;
  wire seg_3_6_sp4_h_r_10_15853;
  wire seg_3_6_sp4_h_r_12_12021;
  wire seg_3_6_sp4_h_r_21_12030;
  wire seg_3_6_sp4_h_r_35_7611;
  wire seg_3_6_sp4_h_r_8_15861;
  wire seg_3_6_sp4_h_r_9_15862;
  wire seg_3_6_sp4_r_v_b_34_15751;
  wire seg_3_6_sp4_v_b_12_11786;
  wire seg_3_6_sp4_v_b_22_11796;
  wire seg_3_6_sp4_v_b_23_11797;
  wire seg_3_6_sp4_v_b_34_11920;
  wire seg_3_6_sp4_v_b_43_12039;
  wire seg_3_6_sp4_v_b_5_11667;
  wire seg_3_6_sp4_v_b_8_11672;
  wire seg_3_6_sp4_v_t_41_12160;
  wire seg_3_6_sp4_v_t_47_12166;
  wire seg_3_7_glb_netwk_0_5;
  wire seg_3_7_glb_netwk_4_9;
  wire seg_3_7_local_g0_2_15882;
  wire seg_3_7_local_g0_3_15883;
  wire seg_3_7_local_g0_4_15884;
  wire seg_3_7_local_g0_5_15885;
  wire seg_3_7_local_g0_6_15886;
  wire seg_3_7_local_g1_0_15888;
  wire seg_3_7_local_g1_1_15889;
  wire seg_3_7_local_g1_2_15890;
  wire seg_3_7_local_g1_3_15891;
  wire seg_3_7_local_g1_4_15892;
  wire seg_3_7_local_g1_6_15894;
  wire seg_3_7_local_g1_7_15895;
  wire seg_3_7_lutff_1_out_12009;
  wire seg_3_7_lutff_4_out_12012;
  wire seg_3_7_lutff_6_out_12014;
  wire seg_3_7_lutff_7_out_12015;
  wire seg_3_7_neigh_op_bnr_1_15717;
  wire seg_3_7_neigh_op_bnr_2_15718;
  wire seg_3_7_neigh_op_bnr_3_15719;
  wire seg_3_7_neigh_op_bnr_5_15721;
  wire seg_3_7_neigh_op_bnr_6_15722;
  wire seg_3_7_sp4_h_l_38_1598;
  wire seg_3_7_sp4_h_r_10_15976;
  wire seg_3_7_sp4_h_r_1_15975;
  wire seg_3_7_sp4_h_r_20_12154;
  wire seg_3_7_sp4_h_r_23_12145;
  wire seg_3_7_sp4_h_r_26_7759;
  wire seg_3_7_sp4_h_r_2_15978;
  wire seg_3_7_sp4_h_r_6_15982;
  wire seg_3_7_sp4_h_r_8_15984;
  wire seg_3_7_sp4_v_b_0_11787;
  wire seg_3_7_sp4_v_b_11_11796;
  wire seg_3_7_sp4_v_b_12_11909;
  wire seg_3_7_sp4_v_b_16_11913;
  wire seg_3_7_sp4_v_b_19_11916;
  wire seg_3_7_sp4_v_b_20_11917;
  wire seg_3_7_sp4_v_b_22_11919;
  wire seg_3_7_sp4_v_b_3_11788;
  wire seg_3_7_sp4_v_b_8_11795;
  wire seg_3_8_glb_netwk_0_5;
  wire seg_3_8_glb_netwk_7_12;
  wire seg_3_8_local_g0_0_16003;
  wire seg_3_8_local_g0_2_16005;
  wire seg_3_8_local_g1_2_16013;
  wire seg_3_8_local_g2_1_16020;
  wire seg_3_8_local_g2_4_16023;
  wire seg_3_8_local_g3_2_16029;
  wire seg_3_8_lutff_4_out_12135;
  wire seg_3_8_neigh_op_tnl_1_7891;
  wire seg_3_8_neigh_op_tnl_4_7894;
  wire seg_3_8_sp4_h_l_36_1805;
  wire seg_3_8_sp4_h_l_44_1814;
  wire seg_3_8_sp4_h_r_16_12273;
  wire seg_3_8_sp4_h_r_18_12275;
  wire seg_3_8_sp4_h_r_20_12277;
  wire seg_3_8_sp4_r_v_b_18_15869;
  wire seg_3_8_sp4_v_b_11_11919;
  wire seg_3_8_sp4_v_b_18_12038;
  wire seg_3_8_sp4_v_b_32_12164;
  wire seg_3_8_sp4_v_b_46_12288;
  wire seg_3_8_sp4_v_b_9_11917;
  wire seg_3_8_sp4_v_t_47_12412;
  wire seg_3_9_local_g0_1_16127;
  wire seg_3_9_local_g0_3_16129;
  wire seg_3_9_local_g0_4_16130;
  wire seg_3_9_local_g0_6_16132;
  wire seg_3_9_local_g0_7_16133;
  wire seg_3_9_local_g1_0_16134;
  wire seg_3_9_local_g1_1_16135;
  wire seg_3_9_local_g1_4_16138;
  wire seg_3_9_local_g1_5_16139;
  wire seg_3_9_local_g1_7_16141;
  wire seg_3_9_local_g2_0_16142;
  wire seg_3_9_local_g2_7_16149;
  wire seg_3_9_local_g3_3_16153;
  wire seg_3_9_local_g3_6_16156;
  wire seg_3_9_lutff_1_out_12255;
  wire seg_3_9_lutff_2_out_12256;
  wire seg_3_9_lutff_3_out_12257;
  wire seg_3_9_lutff_4_out_12258;
  wire seg_3_9_lutff_5_out_12259;
  wire seg_3_9_lutff_6_out_12260;
  wire seg_3_9_lutff_7_out_12261;
  wire seg_3_9_neigh_op_lft_1_7891;
  wire seg_3_9_neigh_op_lft_4_7894;
  wire seg_3_9_neigh_op_lft_5_7895;
  wire seg_3_9_neigh_op_tnl_0_8037;
  wire seg_3_9_neigh_op_tnl_6_8043;
  wire seg_3_9_neigh_op_tnl_7_8044;
  wire seg_3_9_neigh_op_top_0_12377;
  wire seg_3_9_neigh_op_top_1_12378;
  wire seg_3_9_neigh_op_top_3_12380;
  wire seg_3_9_neigh_op_top_4_12381;
  wire seg_3_9_neigh_op_top_7_12384;
  wire seg_3_9_sp4_h_r_11_16223;
  wire seg_3_9_sp4_h_r_3_16225;
  wire seg_3_9_sp4_h_r_5_16227;
  wire seg_3_9_sp4_h_r_6_16228;
  wire seg_3_9_sp4_h_r_9_16231;
  wire seg_3_9_sp4_v_b_15_12158;
  wire seg_3_9_sp4_v_b_43_12408;
  wire seg_3_9_sp4_v_t_36_12524;
  wire seg_3_9_sp4_v_t_43_12531;
  wire seg_3_9_sp4_v_t_46_12534;
  wire seg_4_0_span4_horz_r_0_18923;
  wire seg_4_10_glb_netwk_0_5;
  wire seg_4_10_glb_netwk_4_9;
  wire seg_4_10_local_g2_5_20101;
  wire seg_4_10_local_g3_7_20111;
  wire seg_4_10_neigh_op_bnl_7_12261;
  wire seg_4_10_sp4_h_l_36_2239;
  wire seg_4_10_sp4_h_l_47_2240;
  wire seg_4_10_sp4_h_r_0_20174;
  wire seg_4_10_sp4_h_r_20_16354;
  wire seg_4_10_sp4_h_r_22_16346;
  wire seg_4_10_sp4_h_r_26_12516;
  wire seg_4_10_sp4_h_r_5_20181;
  wire seg_4_10_sp4_r_v_b_47_20197;
  wire seg_4_10_sp4_v_b_24_16233;
  wire seg_4_10_sp4_v_b_28_16237;
  wire seg_4_10_sp4_v_b_32_16241;
  wire seg_4_10_sp4_v_b_34_16243;
  wire seg_4_10_sp4_v_b_37_16356;
  wire seg_4_10_sp4_v_t_41_16483;
  wire seg_4_10_sp4_v_t_42_16484;
  wire seg_4_10_sp4_v_t_44_16486;
  wire seg_4_11_glb_netwk_0_5;
  wire seg_4_11_glb_netwk_4_9;
  wire seg_4_11_local_g0_1_20204;
  wire seg_4_11_local_g0_2_20205;
  wire seg_4_11_local_g0_4_20207;
  wire seg_4_11_local_g1_2_20213;
  wire seg_4_11_local_g1_4_20215;
  wire seg_4_11_local_g2_1_20220;
  wire seg_4_11_local_g3_1_20228;
  wire seg_4_11_local_g3_5_20232;
  wire seg_4_11_sp4_h_l_36_2445;
  wire seg_4_11_sp4_h_l_37_2444;
  wire seg_4_11_sp4_h_l_39_2456;
  wire seg_4_11_sp4_h_l_41_2478;
  wire seg_4_11_sp4_h_l_43_2488;
  wire seg_4_11_sp4_h_l_45_2490;
  wire seg_4_11_sp4_h_l_46_2447;
  wire seg_4_11_sp4_h_l_47_2446;
  wire seg_4_11_sp4_h_r_1_20298;
  wire seg_4_11_sp4_h_r_20_16477;
  wire seg_4_11_sp4_h_r_25_12636;
  wire seg_4_11_sp4_h_r_2_20301;
  wire seg_4_11_sp4_h_r_44_8354;
  wire seg_4_11_sp4_h_r_4_20303;
  wire seg_4_11_sp4_r_v_b_21_20072;
  wire seg_4_11_sp4_r_v_b_25_20186;
  wire seg_4_11_sp4_r_v_b_43_20316;
  wire seg_4_11_sp4_v_b_0_16110;
  wire seg_4_11_sp4_v_b_20_16240;
  wire seg_4_11_sp4_v_b_22_16242;
  wire seg_4_11_sp4_v_b_25_16355;
  wire seg_4_11_sp4_v_b_28_16360;
  wire seg_4_11_sp4_v_b_2_16112;
  wire seg_4_11_sp4_v_b_30_16362;
  wire seg_4_11_sp4_v_b_32_16364;
  wire seg_4_11_sp4_v_b_34_16366;
  wire seg_4_11_sp4_v_b_36_16478;
  wire seg_4_11_sp4_v_b_6_16116;
  wire seg_4_11_sp4_v_b_8_16118;
  wire seg_4_11_sp4_v_t_45_16610;
  wire seg_4_12_glb_netwk_0_5;
  wire seg_4_12_glb_netwk_5_10;
  wire seg_4_12_local_g0_7_20333;
  wire seg_4_12_local_g1_3_20337;
  wire seg_4_12_local_g1_7_20341;
  wire seg_4_12_local_g2_2_20344;
  wire seg_4_12_local_g2_6_20348;
  wire seg_4_12_local_g3_0_20350;
  wire seg_4_12_local_g3_2_20352;
  wire seg_4_12_lutff_2_out_16456;
  wire seg_4_12_neigh_op_tnr_0_20408;
  wire seg_4_12_neigh_op_tnr_2_20410;
  wire seg_4_12_sp4_h_r_10_20422;
  wire seg_4_12_sp4_h_r_15_16593;
  wire seg_4_12_sp4_h_r_18_16598;
  wire seg_4_12_sp4_h_r_24_12758;
  wire seg_4_12_sp4_h_r_2_20424;
  wire seg_4_12_sp4_h_r_34_12760;
  wire seg_4_12_sp4_h_r_4_20426;
  wire seg_4_12_sp4_h_r_6_20428;
  wire seg_4_12_sp4_h_r_8_20430;
  wire seg_4_12_sp4_r_v_b_27_20311;
  wire seg_4_12_sp4_r_v_b_39_20435;
  wire seg_4_12_sp4_v_b_0_16233;
  wire seg_4_12_sp4_v_b_10_16243;
  wire seg_4_12_sp4_v_b_11_16242;
  wire seg_4_12_sp4_v_b_15_16358;
  wire seg_4_12_sp4_v_b_26_16481;
  wire seg_4_12_sp4_v_b_32_16487;
  wire seg_4_12_sp4_v_b_38_16603;
  wire seg_4_12_sp4_v_b_46_16611;
  wire seg_4_12_sp4_v_b_4_16237;
  wire seg_4_12_sp4_v_b_8_16241;
  wire seg_4_13_local_g0_0_20449;
  wire seg_4_13_local_g0_1_20450;
  wire seg_4_13_local_g0_3_20452;
  wire seg_4_13_local_g0_4_20453;
  wire seg_4_13_local_g0_6_20455;
  wire seg_4_13_local_g1_2_20459;
  wire seg_4_13_local_g1_3_20460;
  wire seg_4_13_local_g2_1_20466;
  wire seg_4_13_local_g2_5_20470;
  wire seg_4_13_local_g2_6_20471;
  wire seg_4_13_local_g2_7_20472;
  wire seg_4_13_local_g3_3_20476;
  wire seg_4_13_local_g3_4_20477;
  wire seg_4_13_local_g3_5_20478;
  wire seg_4_13_sp4_h_l_37_2861;
  wire seg_4_13_sp4_h_l_39_2873;
  wire seg_4_13_sp4_h_l_46_2864;
  wire seg_4_13_sp4_h_r_11_20546;
  wire seg_4_13_sp4_h_r_14_16717;
  wire seg_4_13_sp4_h_r_16_16719;
  wire seg_4_13_sp4_h_r_17_16718;
  wire seg_4_13_sp4_h_r_19_16720;
  wire seg_4_13_sp4_h_r_28_12887;
  wire seg_4_13_sp4_h_r_30_12889;
  wire seg_4_13_sp4_h_r_37_8637;
  wire seg_4_13_sp4_h_r_39_8641;
  wire seg_4_13_sp4_h_r_41_8643;
  wire seg_4_13_sp4_h_r_45_8647;
  wire seg_4_13_sp4_h_r_7_20552;
  wire seg_4_13_sp4_r_v_b_19_20316;
  wire seg_4_13_sp4_v_b_10_16366;
  wire seg_4_13_sp4_v_b_11_16365;
  wire seg_4_13_sp4_v_b_12_16478;
  wire seg_4_13_sp4_v_b_3_16357;
  wire seg_4_13_sp4_v_b_4_16360;
  wire seg_4_13_sp4_v_b_5_16359;
  wire seg_4_13_sp4_v_b_6_16362;
  wire seg_4_13_sp4_v_b_8_16364;
  wire seg_4_13_sp4_v_b_9_16363;
  wire seg_4_13_sp4_v_t_41_16852;
  wire seg_4_14_glb_netwk_0_5;
  wire seg_4_14_glb_netwk_4_9;
  wire seg_4_14_local_g1_4_20584;
  wire seg_4_14_local_g2_3_20591;
  wire seg_4_14_local_g2_5_20593;
  wire seg_4_14_local_g3_0_20596;
  wire seg_4_14_local_g3_2_20598;
  wire seg_4_14_local_g3_5_20601;
  wire seg_4_14_local_g3_6_20602;
  wire seg_4_14_lutff_0_out_16700;
  wire seg_4_14_lutff_3_out_16703;
  wire seg_4_14_lutff_4_out_16704;
  wire seg_4_14_lutff_5_out_16705;
  wire seg_4_14_lutff_6_out_16706;
  wire seg_4_14_sp4_h_r_34_13006;
  wire seg_4_14_sp4_h_r_9_20677;
  wire seg_4_14_sp4_r_v_b_3_20311;
  wire seg_4_14_sp4_v_b_14_16603;
  wire seg_4_14_sp4_v_b_27_16726;
  wire seg_4_14_sp4_v_b_2_16481;
  wire seg_4_14_sp4_v_b_32_16733;
  wire seg_4_14_sp4_v_b_45_16856;
  wire seg_4_14_sp4_v_b_5_16482;
  wire seg_4_14_sp4_v_b_8_16487;
  wire seg_4_14_sp4_v_t_36_16970;
  wire seg_4_14_sp4_v_t_43_16977;
  wire seg_4_14_sp4_v_t_46_16980;
  wire seg_4_15_glb_netwk_0_5;
  wire seg_4_15_glb_netwk_4_9;
  wire seg_4_15_local_g0_0_20695;
  wire seg_4_15_local_g2_1_20712;
  wire seg_4_15_local_g2_2_20713;
  wire seg_4_15_local_g2_4_20715;
  wire seg_4_15_local_g2_6_20717;
  wire seg_4_15_local_g3_2_20721;
  wire seg_4_15_local_g3_6_20725;
  wire seg_4_15_local_g3_7_20726;
  wire seg_4_15_lutff_0_out_16823;
  wire seg_4_15_lutff_1_out_16824;
  wire seg_4_15_lutff_2_out_16825;
  wire seg_4_15_lutff_3_out_16826;
  wire seg_4_15_lutff_4_out_16827;
  wire seg_4_15_lutff_5_out_16828;
  wire seg_4_15_lutff_6_out_16829;
  wire seg_4_15_lutff_7_out_16830;
  wire seg_4_15_neigh_op_rgt_4_20658;
  wire seg_4_15_sp4_h_l_45_3344;
  wire seg_4_15_sp4_h_l_47_3300;
  wire seg_4_15_sp4_h_r_34_13129;
  wire seg_4_15_sp4_h_r_38_8936;
  wire seg_4_15_sp4_v_b_0_16602;
  wire seg_4_15_sp4_v_b_11_16611;
  wire seg_4_15_sp4_v_b_34_16858;
  wire seg_4_15_sp4_v_b_4_16606;
  wire seg_4_15_sp4_v_t_37_17094;
  wire seg_4_16_glb_netwk_0_5;
  wire seg_4_16_glb_netwk_4_9;
  wire seg_4_16_local_g0_0_20818;
  wire seg_4_16_local_g0_7_20825;
  wire seg_4_16_local_g1_5_20831;
  wire seg_4_16_local_g2_0_20834;
  wire seg_4_16_local_g2_7_20841;
  wire seg_4_16_local_g3_4_20846;
  wire seg_4_16_lutff_0_out_16946;
  wire seg_4_16_lutff_1_out_16947;
  wire seg_4_16_lutff_4_out_16950;
  wire seg_4_16_lutff_5_out_16951;
  wire seg_4_16_lutff_6_out_16952;
  wire seg_4_16_lutff_7_out_16953;
  wire seg_4_16_sp4_h_l_44_3551;
  wire seg_4_16_sp4_h_r_39_9082;
  wire seg_4_16_sp4_v_b_24_16971;
  wire seg_4_16_sp4_v_t_38_17218;
  wire seg_4_16_sp4_v_t_40_17220;
  wire seg_4_17_glb_netwk_0_5;
  wire seg_4_17_glb_netwk_4_9;
  wire seg_4_17_local_g0_1_20942;
  wire seg_4_17_local_g1_0_20949;
  wire seg_4_17_local_g1_3_20952;
  wire seg_4_17_local_g1_5_20954;
  wire seg_4_17_local_g1_6_20955;
  wire seg_4_17_local_g2_1_20958;
  wire seg_4_17_local_g3_2_20967;
  wire seg_4_17_lutff_1_out_17070;
  wire seg_4_17_lutff_3_out_17072;
  wire seg_4_17_lutff_5_out_17074;
  wire seg_4_17_sp12_h_r_0_21031;
  wire seg_4_17_sp4_h_l_41_3746;
  wire seg_4_17_sp4_h_l_45_3758;
  wire seg_4_17_sp4_h_l_47_3714;
  wire seg_4_17_sp4_h_r_0_21035;
  wire seg_4_17_sp4_h_r_11_21038;
  wire seg_4_17_sp4_h_r_12_17205;
  wire seg_4_17_sp4_h_r_3_21040;
  wire seg_4_17_sp4_h_r_6_21043;
  wire seg_4_17_sp4_h_r_8_21045;
  wire seg_4_17_sp4_h_r_9_21046;
  wire seg_4_17_sp4_r_v_b_31_20930;
  wire seg_4_17_sp4_v_b_0_16848;
  wire seg_4_17_sp4_v_b_1_16847;
  wire seg_4_17_sp4_v_b_25_17093;
  wire seg_4_17_sp4_v_b_34_17104;
  wire seg_4_17_sp4_v_b_3_16849;
  wire seg_4_17_sp4_v_b_9_16855;
  wire seg_4_18_glb_netwk_0_5;
  wire seg_4_18_glb_netwk_4_9;
  wire seg_4_18_local_g0_6_21070;
  wire seg_4_18_local_g1_3_21075;
  wire seg_4_18_local_g1_6_21078;
  wire seg_4_18_local_g3_0_21088;
  wire seg_4_18_local_g3_3_21091;
  wire seg_4_18_sp4_h_l_43_3965;
  wire seg_4_18_sp4_r_v_b_16_20928;
  wire seg_4_18_sp4_r_v_b_19_20931;
  wire seg_4_18_sp4_r_v_b_3_20803;
  wire seg_4_18_sp4_r_v_b_6_20808;
  wire seg_4_18_sp4_v_b_14_17095;
  wire seg_4_18_sp4_v_b_6_16977;
  wire seg_4_19_glb_netwk_0_5;
  wire seg_4_19_glb_netwk_4_9;
  wire seg_4_19_local_g0_5_21192;
  wire seg_4_19_local_g1_1_21196;
  wire seg_4_19_local_g2_2_21205;
  wire seg_4_19_lutff_6_out_17321;
  wire seg_4_19_neigh_op_top_5_17443;
  wire seg_4_19_sp12_v_t_23_21280;
  wire seg_4_19_sp4_h_r_1_21282;
  wire seg_4_19_sp4_h_r_42_9528;
  wire seg_4_19_sp4_v_b_14_17218;
  wire seg_4_19_sp4_v_b_16_17220;
  wire seg_4_19_sp4_v_t_36_17585;
  wire seg_4_19_sp4_v_t_37_17586;
  wire seg_4_1_glb_netwk_0_5;
  wire seg_4_1_glb_netwk_4_9;
  wire seg_4_1_local_g0_2_18935;
  wire seg_4_1_local_g0_3_18936;
  wire seg_4_1_local_g0_7_18940;
  wire seg_4_1_local_g1_1_18942;
  wire seg_4_1_local_g1_2_18943;
  wire seg_4_1_local_g1_3_18944;
  wire seg_4_1_local_g1_4_18945;
  wire seg_4_1_local_g1_5_18946;
  wire seg_4_1_local_g1_7_18948;
  wire seg_4_1_local_g2_0_18949;
  wire seg_4_1_local_g2_2_18951;
  wire seg_4_1_local_g2_3_18952;
  wire seg_4_1_local_g2_5_18954;
  wire seg_4_1_local_g3_3_18960;
  wire seg_4_1_local_g3_6_18963;
  wire seg_4_1_lutff_0_out_15060;
  wire seg_4_1_lutff_2_out_15062;
  wire seg_4_1_lutff_3_out_15063;
  wire seg_4_1_lutff_4_out_15064;
  wire seg_4_1_lutff_5_out_15065;
  wire seg_4_1_lutff_6_out_15066;
  wire seg_4_1_lutff_7_out_15067;
  wire seg_4_1_neigh_op_lft_2_11231;
  wire seg_4_1_neigh_op_lft_3_11232;
  wire seg_4_1_neigh_op_lft_7_11236;
  wire seg_4_1_neigh_op_rgt_3_18894;
  wire seg_4_1_neigh_op_top_2_15190;
  wire seg_4_1_neigh_op_top_3_15191;
  wire seg_4_1_neigh_op_top_7_15195;
  wire seg_4_1_sp4_h_r_5_19038;
  wire seg_4_1_sp4_r_v_b_1_19044;
  wire seg_4_1_sp4_r_v_b_22_19058;
  wire seg_4_1_sp4_r_v_b_39_19076;
  wire seg_4_1_sp4_r_v_b_41_19079;
  wire seg_4_1_sp4_r_v_b_43_19081;
  wire seg_4_1_sp4_v_b_37_15243;
  wire seg_4_1_sp4_v_b_38_15244;
  wire seg_4_1_sp4_v_b_40_15247;
  wire seg_4_1_sp4_v_b_43_15250;
  wire seg_4_20_glb_netwk_0_5;
  wire seg_4_20_glb_netwk_4_9;
  wire seg_4_20_local_g0_5_21315;
  wire seg_4_20_local_g0_7_21317;
  wire seg_4_20_lutff_4_out_17442;
  wire seg_4_20_lutff_5_out_17443;
  wire seg_4_20_sp12_v_b_1_19926;
  wire seg_4_20_sp4_h_l_43_4419;
  wire seg_4_20_sp4_v_b_15_17342;
  wire seg_4_20_sp4_v_b_21_17348;
  wire seg_4_21_sp4_v_b_0_17340;
  wire seg_4_21_sp4_v_b_11_17349;
  wire seg_4_21_sp4_v_b_1_17339;
  wire seg_4_21_sp4_v_b_9_17347;
  wire seg_4_21_sp4_v_t_37_17832;
  wire seg_4_21_sp4_v_t_43_17838;
  wire seg_4_22_glb_netwk_0_5;
  wire seg_4_22_glb_netwk_4_9;
  wire seg_4_22_local_g2_7_21579;
  wire seg_4_22_sp4_h_r_5_21657;
  wire seg_4_22_sp4_v_b_12_17585;
  wire seg_4_22_sp4_v_b_39_17834;
  wire seg_4_23_sp4_h_l_37_5039;
  wire seg_4_25_sp4_h_l_37_5453;
  wire seg_4_25_sp4_h_l_43_5497;
  wire seg_4_25_sp4_h_l_45_5499;
  wire seg_4_2_local_g0_2_19098;
  wire seg_4_2_local_g0_4_19100;
  wire seg_4_2_local_g0_6_19102;
  wire seg_4_2_local_g0_7_19103;
  wire seg_4_2_local_g1_3_19107;
  wire seg_4_2_local_g1_4_19108;
  wire seg_4_2_local_g1_5_19109;
  wire seg_4_2_local_g1_6_19110;
  wire seg_4_2_local_g2_1_19113;
  wire seg_4_2_local_g2_2_19114;
  wire seg_4_2_local_g2_5_19117;
  wire seg_4_2_local_g2_6_19118;
  wire seg_4_2_local_g2_7_19119;
  wire seg_4_2_local_g3_2_19122;
  wire seg_4_2_local_g3_3_19123;
  wire seg_4_2_local_g3_4_19124;
  wire seg_4_2_local_g3_6_19126;
  wire seg_4_2_local_g3_7_19127;
  wire seg_4_2_lutff_1_out_15189;
  wire seg_4_2_lutff_2_out_15190;
  wire seg_4_2_lutff_3_out_15191;
  wire seg_4_2_lutff_4_out_15192;
  wire seg_4_2_lutff_5_out_15193;
  wire seg_4_2_lutff_6_out_15194;
  wire seg_4_2_lutff_7_out_15195;
  wire seg_4_2_neigh_op_bnl_1_11230;
  wire seg_4_2_neigh_op_bnl_2_11231;
  wire seg_4_2_neigh_op_bnl_3_11232;
  wire seg_4_2_neigh_op_bnl_7_11236;
  wire seg_4_2_neigh_op_lft_2_11359;
  wire seg_4_2_neigh_op_lft_4_11361;
  wire seg_4_2_neigh_op_lft_7_11364;
  wire seg_4_2_neigh_op_top_6_15353;
  wire seg_4_2_sp4_h_r_13_15359;
  wire seg_4_2_sp4_h_r_14_15364;
  wire seg_4_2_sp4_h_r_26_11532;
  wire seg_4_2_sp4_r_v_b_13_19060;
  wire seg_4_2_sp4_r_v_b_3_19049;
  wire seg_4_2_sp4_v_b_12_15230;
  wire seg_4_2_sp4_v_b_30_15250;
  wire seg_4_2_sp4_v_b_44_15379;
  wire seg_4_2_sp4_v_b_47_15382;
  wire seg_4_31_span12_vert_0_21280;
  wire seg_4_3_glb_netwk_0_5;
  wire seg_4_3_glb_netwk_4_9;
  wire seg_4_3_local_g0_0_19219;
  wire seg_4_3_local_g0_2_19221;
  wire seg_4_3_local_g0_3_19222;
  wire seg_4_3_local_g0_4_19223;
  wire seg_4_3_local_g0_5_19224;
  wire seg_4_3_local_g0_6_19225;
  wire seg_4_3_local_g1_3_19230;
  wire seg_4_3_local_g1_4_19231;
  wire seg_4_3_local_g1_5_19232;
  wire seg_4_3_local_g1_6_19233;
  wire seg_4_3_local_g1_7_19234;
  wire seg_4_3_local_g2_1_19236;
  wire seg_4_3_local_g2_2_19237;
  wire seg_4_3_local_g2_4_19239;
  wire seg_4_3_local_g2_5_19240;
  wire seg_4_3_local_g2_6_19241;
  wire seg_4_3_local_g2_7_19242;
  wire seg_4_3_local_g3_2_19245;
  wire seg_4_3_local_g3_4_19247;
  wire seg_4_3_local_g3_7_19250;
  wire seg_4_3_lutff_0_out_15347;
  wire seg_4_3_lutff_1_out_15348;
  wire seg_4_3_lutff_2_out_15349;
  wire seg_4_3_lutff_3_out_15350;
  wire seg_4_3_lutff_4_out_15351;
  wire seg_4_3_lutff_5_out_15352;
  wire seg_4_3_lutff_6_out_15353;
  wire seg_4_3_lutff_7_out_15354;
  wire seg_4_3_neigh_op_bnl_6_11363;
  wire seg_4_3_neigh_op_lft_2_11518;
  wire seg_4_3_neigh_op_lft_3_11519;
  wire seg_4_3_neigh_op_lft_4_11520;
  wire seg_4_3_neigh_op_tnl_2_11641;
  wire seg_4_3_neigh_op_top_3_15473;
  wire seg_4_3_neigh_op_top_6_15476;
  wire seg_4_3_sp4_h_l_44_788;
  wire seg_4_3_sp4_h_r_15_15486;
  wire seg_4_3_sp4_h_r_16_15489;
  wire seg_4_3_sp4_h_r_22_15485;
  wire seg_4_3_sp4_h_r_28_11657;
  wire seg_4_3_sp4_h_r_42_7176;
  wire seg_4_3_sp4_r_v_b_13_19074;
  wire seg_4_3_sp4_r_v_b_15_19076;
  wire seg_4_3_sp4_r_v_b_4_19064;
  wire seg_4_3_sp4_v_b_0_15229;
  wire seg_4_3_sp4_v_b_28_15376;
  wire seg_4_3_sp4_v_b_5_15234;
  wire seg_4_3_sp4_v_t_41_15622;
  wire seg_4_3_sp4_v_t_44_15625;
  wire seg_4_4_glb_netwk_0_5;
  wire seg_4_4_glb_netwk_4_9;
  wire seg_4_4_local_g0_4_19346;
  wire seg_4_4_local_g0_6_19348;
  wire seg_4_4_local_g1_0_19350;
  wire seg_4_4_local_g1_2_19352;
  wire seg_4_4_local_g1_3_19353;
  wire seg_4_4_local_g1_4_19354;
  wire seg_4_4_local_g1_6_19356;
  wire seg_4_4_local_g2_2_19360;
  wire seg_4_4_local_g2_3_19361;
  wire seg_4_4_local_g2_4_19362;
  wire seg_4_4_local_g2_7_19365;
  wire seg_4_4_local_g3_5_19371;
  wire seg_4_4_local_g3_7_19373;
  wire seg_4_4_lutff_0_out_15470;
  wire seg_4_4_lutff_3_out_15473;
  wire seg_4_4_lutff_4_out_15474;
  wire seg_4_4_lutff_6_out_15476;
  wire seg_4_4_neigh_op_bot_6_15353;
  wire seg_4_4_neigh_op_lft_2_11641;
  wire seg_4_4_neigh_op_tnl_2_11764;
  wire seg_4_4_sp4_h_l_36_969;
  wire seg_4_4_sp4_h_l_39_980;
  wire seg_4_4_sp4_h_l_47_970;
  wire seg_4_4_sp4_h_r_10_19438;
  wire seg_4_4_sp4_h_r_26_11778;
  wire seg_4_4_sp4_h_r_29_11781;
  wire seg_4_4_sp4_h_r_2_19440;
  wire seg_4_4_sp4_h_r_4_19442;
  wire seg_4_4_sp4_h_r_7_19445;
  wire seg_4_4_sp4_r_v_b_23_19213;
  wire seg_4_4_sp4_r_v_b_28_19330;
  wire seg_4_4_sp4_r_v_b_4_19079;
  wire seg_4_4_sp4_r_v_b_7_19080;
  wire seg_4_4_sp4_v_b_0_15243;
  wire seg_4_4_sp4_v_b_14_15373;
  wire seg_4_4_sp4_v_b_1_15242;
  wire seg_4_4_sp4_v_b_47_15628;
  wire seg_4_4_sp4_v_b_5_15247;
  wire seg_4_4_sp4_v_b_6_15250;
  wire seg_4_4_sp4_v_b_7_15249;
  wire seg_4_4_sp4_v_t_45_15749;
  wire seg_4_5_glb_netwk_0_5;
  wire seg_4_5_glb_netwk_4_9;
  wire seg_4_5_local_g0_5_19470;
  wire seg_4_5_local_g0_6_19471;
  wire seg_4_5_local_g1_0_19473;
  wire seg_4_5_local_g1_1_19474;
  wire seg_4_5_local_g1_5_19478;
  wire seg_4_5_local_g1_6_19479;
  wire seg_4_5_local_g2_0_19481;
  wire seg_4_5_local_g2_2_19483;
  wire seg_4_5_local_g2_4_19485;
  wire seg_4_5_local_g2_7_19488;
  wire seg_4_5_local_g3_3_19492;
  wire seg_4_5_local_g3_4_19493;
  wire seg_4_5_local_g3_5_19494;
  wire seg_4_5_local_g3_6_19495;
  wire seg_4_5_local_g3_7_19496;
  wire seg_4_5_lutff_0_out_15593;
  wire seg_4_5_lutff_3_out_15596;
  wire seg_4_5_lutff_4_out_15597;
  wire seg_4_5_lutff_5_out_15598;
  wire seg_4_5_lutff_6_out_15599;
  wire seg_4_5_lutff_7_out_15600;
  wire seg_4_5_neigh_op_bnl_0_11639;
  wire seg_4_5_neigh_op_bnr_6_19307;
  wire seg_4_5_neigh_op_rgt_7_19431;
  wire seg_4_5_sp4_h_l_37_1178;
  wire seg_4_5_sp4_h_l_43_1222;
  wire seg_4_5_sp4_h_l_44_1225;
  wire seg_4_5_sp4_h_r_10_19561;
  wire seg_4_5_sp4_h_r_12_15729;
  wire seg_4_5_sp4_h_r_18_15737;
  wire seg_4_5_sp4_h_r_1_19560;
  wire seg_4_5_sp4_h_r_20_15739;
  wire seg_4_5_sp4_h_r_28_11903;
  wire seg_4_5_sp4_h_r_31_11906;
  wire seg_4_5_sp4_h_r_34_11899;
  wire seg_4_5_sp4_h_r_4_19565;
  wire seg_4_5_sp4_r_v_b_36_19571;
  wire seg_4_5_sp4_r_v_b_46_19581;
  wire seg_4_5_sp4_v_b_28_15622;
  wire seg_4_5_sp4_v_b_35_15627;
  wire seg_4_5_sp4_v_b_37_15741;
  wire seg_4_5_sp4_v_b_42_15746;
  wire seg_4_5_sp4_v_b_44_15748;
  wire seg_4_5_sp4_v_b_5_15375;
  wire seg_4_5_sp4_v_t_36_15863;
  wire seg_4_5_sp4_v_t_47_15874;
  wire seg_4_6_glb_netwk_0_5;
  wire seg_4_6_glb_netwk_3_8;
  wire seg_4_6_local_g0_0_19588;
  wire seg_4_6_local_g0_2_19590;
  wire seg_4_6_local_g0_3_19591;
  wire seg_4_6_local_g0_4_19592;
  wire seg_4_6_local_g0_7_19595;
  wire seg_4_6_local_g1_0_19596;
  wire seg_4_6_local_g1_3_19599;
  wire seg_4_6_local_g1_6_19602;
  wire seg_4_6_local_g1_7_19603;
  wire seg_4_6_local_g2_0_19604;
  wire seg_4_6_local_g3_0_19612;
  wire seg_4_6_local_g3_3_19615;
  wire seg_4_6_lutff_0_out_15716;
  wire seg_4_6_lutff_1_out_15717;
  wire seg_4_6_lutff_2_out_15718;
  wire seg_4_6_lutff_3_out_15719;
  wire seg_4_6_lutff_5_out_15721;
  wire seg_4_6_lutff_6_out_15722;
  wire seg_4_6_lutff_7_out_15723;
  wire seg_4_6_neigh_op_lft_0_11885;
  wire seg_4_6_sp4_h_l_37_1384;
  wire seg_4_6_sp4_h_l_41_1418;
  wire seg_4_6_sp4_h_l_42_1429;
  wire seg_4_6_sp4_h_l_47_1386;
  wire seg_4_6_sp4_h_r_10_19684;
  wire seg_4_6_sp4_h_r_20_15862;
  wire seg_4_6_sp4_h_r_32_12030;
  wire seg_4_6_sp4_h_r_3_19687;
  wire seg_4_6_sp4_h_r_5_19689;
  wire seg_4_6_sp4_h_r_7_19691;
  wire seg_4_6_sp4_h_r_9_19693;
  wire seg_4_6_sp4_r_v_b_16_19452;
  wire seg_4_6_sp4_r_v_b_19_19455;
  wire seg_4_6_sp4_r_v_b_24_19572;
  wire seg_4_6_sp4_r_v_b_32_19580;
  wire seg_4_6_sp4_r_v_b_41_19699;
  wire seg_4_6_sp4_r_v_b_6_19332;
  wire seg_4_6_sp4_v_t_38_15988;
  wire seg_4_6_sp4_v_t_40_15990;
  wire seg_4_6_sp4_v_t_42_15992;
  wire seg_4_7_glb_netwk_0_5;
  wire seg_4_7_glb_netwk_3_8;
  wire seg_4_7_local_g0_1_19712;
  wire seg_4_7_local_g0_4_19715;
  wire seg_4_7_local_g0_7_19718;
  wire seg_4_7_local_g1_1_19720;
  wire seg_4_7_local_g1_2_19721;
  wire seg_4_7_local_g1_5_19724;
  wire seg_4_7_local_g1_6_19725;
  wire seg_4_7_local_g1_7_19726;
  wire seg_4_7_local_g2_2_19729;
  wire seg_4_7_local_g2_4_19731;
  wire seg_4_7_local_g2_5_19732;
  wire seg_4_7_local_g2_7_19734;
  wire seg_4_7_local_g3_0_19735;
  wire seg_4_7_local_g3_1_19736;
  wire seg_4_7_local_g3_2_19737;
  wire seg_4_7_local_g3_3_19738;
  wire seg_4_7_local_g3_5_19740;
  wire seg_4_7_local_g3_7_19742;
  wire seg_4_7_lutff_1_out_15840;
  wire seg_4_7_lutff_3_out_15842;
  wire seg_4_7_lutff_5_out_15844;
  wire seg_4_7_lutff_6_out_15845;
  wire seg_4_7_lutff_7_out_15846;
  wire seg_4_7_neigh_op_bnl_5_11890;
  wire seg_4_7_neigh_op_bnl_7_11892;
  wire seg_4_7_neigh_op_rgt_3_19673;
  wire seg_4_7_sp4_h_l_39_1604;
  wire seg_4_7_sp4_h_l_43_1636;
  wire seg_4_7_sp4_h_l_46_1595;
  wire seg_4_7_sp4_h_l_47_1594;
  wire seg_4_7_sp4_h_r_0_19805;
  wire seg_4_7_sp4_h_r_23_15976;
  wire seg_4_7_sp4_h_r_4_19811;
  wire seg_4_7_sp4_h_r_8_19815;
  wire seg_4_7_sp4_r_v_b_10_19459;
  wire seg_4_7_sp4_r_v_b_16_19575;
  wire seg_4_7_sp4_r_v_b_17_19576;
  wire seg_4_7_sp4_r_v_b_18_19577;
  wire seg_4_7_sp4_r_v_b_23_19582;
  wire seg_4_7_sp4_r_v_b_29_19698;
  wire seg_4_7_sp4_r_v_b_36_19817;
  wire seg_4_7_sp4_r_v_b_37_19818;
  wire seg_4_7_sp4_r_v_b_9_19456;
  wire seg_4_7_sp4_v_b_17_15745;
  wire seg_4_7_sp4_v_b_18_15746;
  wire seg_4_7_sp4_v_b_20_15748;
  wire seg_4_7_sp4_v_t_36_16109;
  wire seg_4_7_sp4_v_t_38_16111;
  wire seg_4_7_sp4_v_t_42_16115;
  wire seg_4_7_sp4_v_t_43_16116;
  wire seg_4_7_sp4_v_t_45_16118;
  wire seg_4_7_sp4_v_t_46_16119;
  wire seg_4_8_glb_netwk_0_5;
  wire seg_4_8_glb_netwk_4_9;
  wire seg_4_8_local_g0_4_19838;
  wire seg_4_8_local_g1_6_19848;
  wire seg_4_8_local_g2_2_19852;
  wire seg_4_8_local_g2_4_19854;
  wire seg_4_8_local_g2_6_19856;
  wire seg_4_8_local_g3_1_19859;
  wire seg_4_8_local_g3_3_19861;
  wire seg_4_8_local_g3_5_19863;
  wire seg_4_8_local_g3_7_19865;
  wire seg_4_8_neigh_op_lft_4_12135;
  wire seg_4_8_neigh_op_tnl_1_12255;
  wire seg_4_8_neigh_op_tnl_2_12256;
  wire seg_4_8_neigh_op_tnl_3_12257;
  wire seg_4_8_neigh_op_tnl_4_12258;
  wire seg_4_8_neigh_op_tnl_5_12259;
  wire seg_4_8_neigh_op_tnl_6_12260;
  wire seg_4_8_neigh_op_tnl_7_12261;
  wire seg_4_8_sp12_h_r_1_19925;
  wire seg_4_8_sp12_v_b_23_19804;
  wire seg_4_8_sp4_h_l_37_1801;
  wire seg_4_8_sp4_h_r_10_19930;
  wire seg_4_8_sp4_h_r_11_19931;
  wire seg_4_8_sp4_h_r_2_19932;
  wire seg_4_8_sp4_h_r_5_19935;
  wire seg_4_8_sp4_r_v_b_47_19951;
  wire seg_4_8_sp4_v_b_14_15865;
  wire seg_4_8_sp4_v_b_1_15740;
  wire seg_4_8_sp4_v_t_40_16236;
  wire seg_4_9_glb_netwk_0_5;
  wire seg_4_9_glb_netwk_4_9;
  wire seg_4_9_local_g0_3_19960;
  wire seg_4_9_local_g1_7_19972;
  wire seg_4_9_neigh_op_lft_7_12261;
  wire seg_4_9_sp4_h_r_0_20051;
  wire seg_4_9_sp4_h_r_10_20053;
  wire seg_4_9_sp4_h_r_11_20054;
  wire seg_4_9_sp4_h_r_14_16225;
  wire seg_4_9_sp4_h_r_20_16231;
  wire seg_4_9_sp4_h_r_22_16223;
  wire seg_4_9_sp4_h_r_24_12389;
  wire seg_4_9_sp4_h_r_32_12399;
  wire seg_4_9_sp4_h_r_5_20058;
  wire seg_4_9_sp4_h_r_6_20059;
  wire seg_4_9_sp4_h_r_8_20061;
  wire seg_4_9_sp4_h_r_9_20062;
  wire seg_4_9_sp4_r_v_b_27_19942;
  wire seg_4_9_sp4_r_v_b_29_19944;
  wire seg_4_9_sp4_r_v_b_35_19950;
  wire seg_4_9_sp4_v_b_3_15865;
  wire seg_4_9_sp4_v_b_5_15867;
  wire seg_4_9_sp4_v_t_37_16356;
  wire seg_4_9_sp4_v_t_42_16361;
  wire seg_4_9_sp4_v_t_45_16364;
  wire seg_5_0_local_g1_7_22721;
  wire seg_5_0_logic_op_top_7_18898;
  wire seg_5_0_span4_horz_r_2_22756;
  wire seg_5_10_glb_netwk_0_5;
  wire seg_5_10_glb_netwk_7_12;
  wire seg_5_10_local_g0_3_23914;
  wire seg_5_10_local_g0_5_23916;
  wire seg_5_10_local_g0_7_23918;
  wire seg_5_10_local_g1_1_23920;
  wire seg_5_10_local_g2_2_23929;
  wire seg_5_10_local_g2_6_23933;
  wire seg_5_10_local_g3_2_23937;
  wire seg_5_10_local_g3_4_23939;
  wire seg_5_10_sp12_v_b_12_23266;
  wire seg_5_10_sp12_v_b_19_23635;
  wire seg_5_10_sp12_v_b_4_22746;
  wire seg_5_10_sp4_h_l_36_8197;
  wire seg_5_10_sp4_h_l_37_8196;
  wire seg_5_10_sp4_h_l_41_8202;
  wire seg_5_10_sp4_h_l_43_8204;
  wire seg_5_10_sp4_h_r_10_24007;
  wire seg_5_10_sp4_h_r_16_20181;
  wire seg_5_10_sp4_h_r_1_24006;
  wire seg_5_10_sp4_h_r_30_16351;
  wire seg_5_10_sp4_h_r_34_16345;
  wire seg_5_10_sp4_h_r_5_24012;
  wire seg_5_10_sp4_h_r_7_24014;
  wire seg_5_10_sp4_h_r_9_24016;
  wire seg_5_10_sp4_r_v_b_15_23774;
  wire seg_5_10_sp4_r_v_b_19_23778;
  wire seg_5_10_sp4_r_v_b_39_24020;
  wire seg_5_10_sp4_v_b_19_19947;
  wire seg_5_10_sp4_v_b_20_19948;
  wire seg_5_10_sp4_v_b_26_20066;
  wire seg_5_10_sp4_v_b_40_20190;
  wire seg_5_10_sp4_v_t_37_20310;
  wire seg_5_10_sp4_v_t_39_20312;
  wire seg_5_10_sp4_v_t_40_20313;
  wire seg_5_10_sp4_v_t_42_20315;
  wire seg_5_10_sp4_v_t_44_20317;
  wire seg_5_10_sp4_v_t_46_20319;
  wire seg_5_11_glb_netwk_0_5;
  wire seg_5_11_glb_netwk_4_9;
  wire seg_5_11_local_g1_0_24042;
  wire seg_5_11_local_g1_7_24049;
  wire seg_5_11_local_g2_0_24050;
  wire seg_5_11_local_g2_2_24052;
  wire seg_5_11_local_g2_4_24054;
  wire seg_5_11_local_g3_0_24058;
  wire seg_5_11_local_g3_2_24060;
  wire seg_5_11_local_g3_4_24062;
  wire seg_5_11_neigh_op_rgt_0_23993;
  wire seg_5_11_neigh_op_rgt_2_23995;
  wire seg_5_11_neigh_op_rgt_4_23997;
  wire seg_5_11_neigh_op_tnr_0_24116;
  wire seg_5_11_neigh_op_tnr_4_24120;
  wire seg_5_11_sp4_h_l_39_8347;
  wire seg_5_11_sp4_h_l_42_8352;
  wire seg_5_11_sp4_h_l_43_8351;
  wire seg_5_11_sp4_h_r_0_24128;
  wire seg_5_11_sp4_h_r_18_20306;
  wire seg_5_11_sp4_h_r_23_20299;
  wire seg_5_11_sp4_h_r_32_16476;
  wire seg_5_11_sp4_h_r_6_24136;
  wire seg_5_11_sp4_r_v_b_10_23782;
  wire seg_5_11_sp4_v_b_0_19941;
  wire seg_5_11_sp4_v_b_10_19951;
  wire seg_5_11_sp4_v_b_11_19950;
  wire seg_5_11_sp4_v_b_24_20187;
  wire seg_5_11_sp4_v_b_26_20189;
  wire seg_5_11_sp4_v_b_28_20191;
  wire seg_5_11_sp4_v_b_32_20195;
  wire seg_5_11_sp4_v_b_36_20309;
  wire seg_5_11_sp4_v_b_3_19942;
  wire seg_5_11_sp4_v_b_46_20319;
  wire seg_5_11_sp4_v_b_4_19945;
  wire seg_5_11_sp4_v_b_5_19944;
  wire seg_5_11_sp4_v_b_9_19948;
  wire seg_5_12_glb_netwk_0_5;
  wire seg_5_12_glb_netwk_4_9;
  wire seg_5_12_local_g0_4_24161;
  wire seg_5_12_local_g0_7_24164;
  wire seg_5_12_local_g1_5_24170;
  wire seg_5_12_local_g2_0_24173;
  wire seg_5_12_local_g2_2_24175;
  wire seg_5_12_local_g2_4_24177;
  wire seg_5_12_local_g3_1_24182;
  wire seg_5_12_local_g3_3_24184;
  wire seg_5_12_lutff_2_out_20287;
  wire seg_5_12_lutff_4_out_20289;
  wire seg_5_12_neigh_op_bnr_5_23998;
  wire seg_5_12_neigh_op_top_4_20412;
  wire seg_5_12_neigh_op_top_7_20415;
  wire seg_5_12_sp12_v_b_0_22746;
  wire seg_5_12_sp4_h_r_18_20429;
  wire seg_5_12_sp4_h_r_1_24252;
  wire seg_5_12_sp4_h_r_22_20423;
  wire seg_5_12_sp4_h_r_24_16589;
  wire seg_5_12_sp4_h_r_28_16595;
  wire seg_5_12_sp4_h_r_32_16599;
  wire seg_5_12_sp4_h_r_34_16591;
  wire seg_5_12_sp4_h_r_35_16592;
  wire seg_5_12_sp4_h_r_3_24256;
  wire seg_5_12_sp4_h_r_46_12761;
  wire seg_5_12_sp4_h_r_6_24259;
  wire seg_5_12_sp4_r_v_b_19_24024;
  wire seg_5_12_sp4_r_v_b_31_24146;
  wire seg_5_12_sp4_r_v_b_33_24148;
  wire seg_5_12_sp4_v_b_11_20073;
  wire seg_5_12_sp4_v_b_1_20063;
  wire seg_5_12_sp4_v_b_26_20312;
  wire seg_5_12_sp4_v_b_2_20066;
  wire seg_5_12_sp4_v_b_3_20065;
  wire seg_5_12_sp4_v_b_41_20437;
  wire seg_5_12_sp4_v_b_5_20067;
  wire seg_5_12_sp4_v_b_6_20070;
  wire seg_5_12_sp4_v_b_7_20069;
  wire seg_5_12_sp4_v_b_9_20071;
  wire seg_5_12_sp4_v_t_41_20560;
  wire seg_5_12_sp4_v_t_47_20566;
  wire seg_5_13_glb_netwk_0_5;
  wire seg_5_13_glb_netwk_4_9;
  wire seg_5_13_local_g0_3_24283;
  wire seg_5_13_local_g0_6_24286;
  wire seg_5_13_local_g1_5_24293;
  wire seg_5_13_local_g2_0_24296;
  wire seg_5_13_local_g2_2_24298;
  wire seg_5_13_local_g2_4_24300;
  wire seg_5_13_local_g3_2_24306;
  wire seg_5_13_local_g3_6_24310;
  wire seg_5_13_lutff_0_out_20408;
  wire seg_5_13_lutff_2_out_20410;
  wire seg_5_13_lutff_3_out_20411;
  wire seg_5_13_lutff_4_out_20412;
  wire seg_5_13_lutff_5_out_20413;
  wire seg_5_13_lutff_6_out_20414;
  wire seg_5_13_lutff_7_out_20415;
  wire seg_5_13_sp12_v_b_0_22861;
  wire seg_5_13_sp4_h_l_46_8640;
  wire seg_5_13_sp4_h_l_47_8639;
  wire seg_5_13_sp4_h_r_18_20552;
  wire seg_5_13_sp4_h_r_26_16716;
  wire seg_5_13_sp4_h_r_2_24378;
  wire seg_5_13_sp4_h_r_32_16722;
  wire seg_5_13_sp4_h_r_34_16714;
  wire seg_5_13_sp4_h_r_44_12892;
  wire seg_5_13_sp4_h_r_46_12884;
  wire seg_5_13_sp4_r_v_b_17_24145;
  wire seg_5_13_sp4_r_v_b_19_24147;
  wire seg_5_13_sp4_v_b_0_20187;
  wire seg_5_13_sp4_v_b_10_20197;
  wire seg_5_13_sp4_v_b_16_20313;
  wire seg_5_13_sp4_v_b_1_20186;
  wire seg_5_13_sp4_v_b_20_20317;
  wire seg_5_13_sp4_v_b_2_20189;
  wire seg_5_13_sp4_v_b_34_20443;
  wire seg_5_13_sp4_v_b_3_20188;
  wire seg_5_13_sp4_v_b_4_20191;
  wire seg_5_13_sp4_v_b_5_20190;
  wire seg_5_13_sp4_v_b_6_20193;
  wire seg_5_13_sp4_v_b_7_20192;
  wire seg_5_13_sp4_v_b_8_20195;
  wire seg_5_13_sp4_v_b_9_20194;
  wire seg_5_14_glb_netwk_0_5;
  wire seg_5_14_glb_netwk_4_9;
  wire seg_5_14_local_g1_5_24416;
  wire seg_5_14_local_g2_2_24421;
  wire seg_5_14_local_g2_4_24423;
  wire seg_5_14_local_g3_1_24428;
  wire seg_5_14_local_g3_4_24431;
  wire seg_5_14_local_g3_5_24432;
  wire seg_5_14_lutff_1_out_20532;
  wire seg_5_14_lutff_2_out_20533;
  wire seg_5_14_lutff_4_out_20535;
  wire seg_5_14_lutff_5_out_20536;
  wire seg_5_14_sp4_h_l_36_8785;
  wire seg_5_14_sp4_h_r_9_24508;
  wire seg_5_14_sp4_r_v_b_17_24268;
  wire seg_5_14_sp4_r_v_b_20_24271;
  wire seg_5_14_sp4_r_v_b_31_24392;
  wire seg_5_14_sp4_v_b_10_20320;
  wire seg_5_14_sp4_v_b_11_20319;
  wire seg_5_14_sp4_v_b_13_20433;
  wire seg_5_14_sp4_v_b_1_20309;
  wire seg_5_14_sp4_v_b_2_20312;
  wire seg_5_14_sp4_v_t_41_20806;
  wire seg_5_14_sp4_v_t_42_20807;
  wire seg_5_15_glb_netwk_0_5;
  wire seg_5_15_glb_netwk_4_9;
  wire seg_5_15_local_g0_7_24533;
  wire seg_5_15_local_g1_1_24535;
  wire seg_5_15_local_g1_4_24538;
  wire seg_5_15_local_g2_6_24548;
  wire seg_5_15_local_g3_1_24551;
  wire seg_5_15_local_g3_3_24553;
  wire seg_5_15_local_g3_7_24557;
  wire seg_5_15_lutff_1_out_20655;
  wire seg_5_15_lutff_3_out_20657;
  wire seg_5_15_lutff_4_out_20658;
  wire seg_5_15_lutff_6_out_20660;
  wire seg_5_15_lutff_7_out_20661;
  wire seg_5_15_sp4_h_l_41_8937;
  wire seg_5_15_sp4_h_l_47_8933;
  wire seg_5_15_sp4_h_r_0_24620;
  wire seg_5_15_sp4_h_r_1_24621;
  wire seg_5_15_sp4_h_r_4_24626;
  wire seg_5_15_sp4_h_r_7_24629;
  wire seg_5_15_sp4_r_v_b_43_24639;
  wire seg_5_15_sp4_v_b_10_20443;
  wire seg_5_15_sp4_v_b_2_20435;
  wire seg_5_15_sp4_v_b_4_20437;
  wire seg_5_15_sp4_v_b_5_20436;
  wire seg_5_15_sp4_v_t_42_20930;
  wire seg_5_16_glb_netwk_0_5;
  wire seg_5_16_glb_netwk_4_9;
  wire seg_5_16_local_g0_0_24649;
  wire seg_5_16_local_g0_2_24651;
  wire seg_5_16_local_g0_4_24653;
  wire seg_5_16_local_g0_5_24654;
  wire seg_5_16_local_g0_7_24656;
  wire seg_5_16_local_g1_0_24657;
  wire seg_5_16_local_g1_1_24658;
  wire seg_5_16_local_g1_2_24659;
  wire seg_5_16_local_g1_3_24660;
  wire seg_5_16_local_g1_4_24661;
  wire seg_5_16_local_g1_5_24662;
  wire seg_5_16_local_g2_0_24665;
  wire seg_5_16_local_g3_2_24675;
  wire seg_5_16_local_g3_3_24676;
  wire seg_5_16_local_g3_7_24680;
  wire seg_5_16_sp12_v_b_0_23266;
  wire seg_5_16_sp12_v_b_3_23389;
  wire seg_5_16_sp4_h_l_41_9084;
  wire seg_5_16_sp4_h_r_18_20921;
  wire seg_5_16_sp4_r_v_b_15_24512;
  wire seg_5_16_sp4_r_v_b_18_24515;
  wire seg_5_16_sp4_r_v_b_23_24520;
  wire seg_5_16_sp4_r_v_b_27_24634;
  wire seg_5_16_sp4_r_v_b_2_24389;
  wire seg_5_16_sp4_r_v_b_4_24391;
  wire seg_5_16_sp4_r_v_b_5_24390;
  wire seg_5_16_sp4_v_b_0_20556;
  wire seg_5_16_sp4_v_b_10_20566;
  wire seg_5_16_sp4_v_b_13_20679;
  wire seg_5_16_sp4_v_b_16_20682;
  wire seg_5_16_sp4_v_b_1_20555;
  wire seg_5_16_sp4_v_b_20_20686;
  wire seg_5_16_sp4_v_b_23_20689;
  wire seg_5_16_sp4_v_b_28_20806;
  wire seg_5_16_sp4_v_b_3_20557;
  wire seg_5_16_sp4_v_b_4_20560;
  wire seg_5_17_glb_netwk_0_5;
  wire seg_5_17_glb_netwk_4_9;
  wire seg_5_17_local_g0_0_24772;
  wire seg_5_17_local_g0_1_24773;
  wire seg_5_17_local_g1_0_24780;
  wire seg_5_17_local_g1_3_24783;
  wire seg_5_17_local_g2_4_24792;
  wire seg_5_17_lutff_1_out_20901;
  wire seg_5_17_sp4_h_r_0_24866;
  wire seg_5_17_sp4_h_r_2_24870;
  wire seg_5_17_sp4_h_r_34_17206;
  wire seg_5_17_sp4_r_v_b_0_24510;
  wire seg_5_17_sp4_r_v_b_12_24632;
  wire seg_5_17_sp4_v_b_2_20681;
  wire seg_5_17_sp4_v_b_3_20680;
  wire seg_5_17_sp4_v_b_4_20683;
  wire seg_5_17_sp4_v_b_7_20684;
  wire seg_5_17_sp4_v_b_8_20687;
  wire seg_5_18_glb_netwk_0_5;
  wire seg_5_18_glb_netwk_5_10;
  wire seg_5_18_local_g0_0_24895;
  wire seg_5_18_local_g0_4_24899;
  wire seg_5_18_local_g3_6_24925;
  wire seg_5_18_neigh_op_tnl_6_17321;
  wire seg_5_18_neigh_op_top_0_21146;
  wire seg_5_18_sp4_h_r_22_21161;
  wire seg_5_18_sp4_h_r_24_17327;
  wire seg_5_18_sp4_h_r_8_24999;
  wire seg_5_18_sp4_r_v_b_3_24634;
  wire seg_5_18_sp4_v_b_12_20924;
  wire seg_5_18_sp4_v_b_1_20801;
  wire seg_5_18_sp4_v_b_2_20804;
  wire seg_5_18_sp4_v_t_42_21299;
  wire seg_5_19_glb_netwk_0_5;
  wire seg_5_19_glb_netwk_4_9;
  wire seg_5_19_local_g0_6_25024;
  wire seg_5_19_local_g2_4_25038;
  wire seg_5_19_lutff_0_out_21146;
  wire seg_5_19_neigh_op_tnl_4_17442;
  wire seg_5_19_sp12_v_t_23_25111;
  wire seg_5_19_sp4_h_l_38_9524;
  wire seg_5_19_sp4_h_l_40_9526;
  wire seg_5_19_sp4_h_l_41_9525;
  wire seg_5_19_sp4_h_l_44_9530;
  wire seg_5_19_sp4_h_r_24_17450;
  wire seg_5_19_sp4_h_r_6_25120;
  wire seg_5_1_glb_netwk_0_5;
  wire seg_5_1_glb_netwk_4_9;
  wire seg_5_1_local_g2_5_22785;
  wire seg_5_1_local_g3_2_22790;
  wire seg_5_1_local_g3_3_22791;
  wire seg_5_1_lutff_3_out_18894;
  wire seg_5_1_lutff_7_out_18898;
  wire seg_5_1_sp4_h_r_7_22871;
  wire seg_5_1_sp4_r_v_b_13_22879;
  wire seg_5_1_sp4_v_b_42_19080;
  wire seg_5_1_sp4_v_t_47_19213;
  wire seg_5_21_sp4_v_b_3_21172;
  wire seg_5_21_sp4_v_b_5_21174;
  wire seg_5_21_sp4_v_b_7_21176;
  wire seg_5_22_sp4_v_t_41_21790;
  wire seg_5_26_sp4_v_t_36_22277;
  wire seg_5_2_glb_netwk_0_5;
  wire seg_5_2_glb_netwk_3_8;
  wire seg_5_2_local_g2_1_22944;
  wire seg_5_2_local_g3_4_22955;
  wire seg_5_2_lutff_5_out_19024;
  wire seg_5_2_sp12_v_b_11_22734;
  wire seg_5_2_sp12_v_b_20_22746;
  wire seg_5_2_sp4_h_l_46_7023;
  wire seg_5_2_sp4_h_r_10_23023;
  wire seg_5_2_sp4_r_v_b_19_22898;
  wire seg_5_2_sp4_v_b_33_19082;
  wire seg_5_2_sp4_v_t_36_19325;
  wire seg_5_30_sp4_v_t_40_26489;
  wire seg_5_31_span12_vert_0_25111;
  wire seg_5_31_span4_vert_40_26489;
  wire seg_5_3_glb_netwk_0_5;
  wire seg_5_3_local_g0_5_23055;
  wire seg_5_3_local_g0_6_23056;
  wire seg_5_3_local_g1_3_23061;
  wire seg_5_3_local_g1_5_23063;
  wire seg_5_3_local_g2_3_23069;
  wire seg_5_3_local_g2_5_23071;
  wire seg_5_3_local_g3_3_23077;
  wire seg_5_3_local_g3_4_23078;
  wire seg_5_3_lutff_2_out_19180;
  wire seg_5_3_lutff_5_out_19183;
  wire seg_5_3_neigh_op_bot_5_19024;
  wire seg_5_3_sp12_v_b_19_22746;
  wire seg_5_3_sp12_v_b_20_22861;
  wire seg_5_3_sp4_h_l_42_7176;
  wire seg_5_3_sp4_h_l_45_7177;
  wire seg_5_3_sp4_h_l_47_7169;
  wire seg_5_3_sp4_h_r_0_23144;
  wire seg_5_3_sp4_h_r_11_23147;
  wire seg_5_3_sp4_h_r_22_19316;
  wire seg_5_3_sp4_h_r_4_23150;
  wire seg_5_3_sp4_h_r_5_23151;
  wire seg_5_3_sp4_r_v_b_19_22912;
  wire seg_5_3_sp4_v_b_21_19083;
  wire seg_5_3_sp4_v_b_30_19209;
  wire seg_5_3_sp4_v_b_8_19069;
  wire seg_5_3_sp4_v_t_43_19455;
  wire seg_5_3_sp4_v_t_44_19456;
  wire seg_5_3_sp4_v_t_45_19457;
  wire seg_5_3_sp4_v_t_46_19458;
  wire seg_5_4_glb_netwk_0_5;
  wire seg_5_4_glb_netwk_4_9;
  wire seg_5_4_local_g0_4_23177;
  wire seg_5_4_local_g0_6_23179;
  wire seg_5_4_local_g1_5_23186;
  wire seg_5_4_local_g1_7_23188;
  wire seg_5_4_local_g2_0_23189;
  wire seg_5_4_local_g2_1_23190;
  wire seg_5_4_local_g3_0_23197;
  wire seg_5_4_local_g3_1_23198;
  wire seg_5_4_local_g3_7_23204;
  wire seg_5_4_lutff_6_out_19307;
  wire seg_5_4_neigh_op_bnr_4_23013;
  wire seg_5_4_neigh_op_bnr_5_23014;
  wire seg_5_4_neigh_op_bnr_6_23015;
  wire seg_5_4_neigh_op_bnr_7_23016;
  wire seg_5_4_neigh_op_rgt_0_23132;
  wire seg_5_4_neigh_op_rgt_1_23133;
  wire seg_5_4_neigh_op_tnl_7_15600;
  wire seg_5_4_sp4_h_l_37_7314;
  wire seg_5_4_sp4_h_r_11_23270;
  wire seg_5_4_sp4_h_r_14_19441;
  wire seg_5_4_sp4_h_r_4_23273;
  wire seg_5_4_sp4_r_v_b_17_23038;
  wire seg_5_4_sp4_r_v_b_43_23286;
  wire seg_5_4_sp4_r_v_b_45_23288;
  wire seg_5_4_sp4_v_b_24_19326;
  wire seg_5_4_sp4_v_b_32_19334;
  wire seg_5_4_sp4_v_b_34_19336;
  wire seg_5_4_sp4_v_b_36_19448;
  wire seg_5_4_sp4_v_b_38_19450;
  wire seg_5_4_sp4_v_b_40_19452;
  wire seg_5_4_sp4_v_b_6_19081;
  wire seg_5_4_sp4_v_t_37_19572;
  wire seg_5_4_sp4_v_t_43_19578;
  wire seg_5_5_glb_netwk_0_5;
  wire seg_5_5_glb_netwk_4_9;
  wire seg_5_5_local_g0_3_23299;
  wire seg_5_5_local_g0_5_23301;
  wire seg_5_5_local_g1_1_23305;
  wire seg_5_5_local_g1_2_23306;
  wire seg_5_5_local_g1_3_23307;
  wire seg_5_5_local_g1_4_23308;
  wire seg_5_5_local_g1_6_23310;
  wire seg_5_5_local_g3_7_23327;
  wire seg_5_5_lutff_7_out_19431;
  wire seg_5_5_neigh_op_lft_3_15596;
  wire seg_5_5_neigh_op_top_1_19548;
  wire seg_5_5_neigh_op_top_2_19549;
  wire seg_5_5_neigh_op_top_3_19550;
  wire seg_5_5_neigh_op_top_4_19551;
  wire seg_5_5_neigh_op_top_5_19552;
  wire seg_5_5_neigh_op_top_6_19553;
  wire seg_5_5_sp4_h_l_39_7465;
  wire seg_5_5_sp4_h_r_0_23390;
  wire seg_5_5_sp4_h_r_10_23392;
  wire seg_5_5_sp4_h_r_1_23391;
  wire seg_5_5_sp4_h_r_2_23394;
  wire seg_5_5_sp4_h_r_34_15730;
  wire seg_5_5_sp4_h_r_36_11898;
  wire seg_5_5_sp4_h_r_38_11902;
  wire seg_5_5_sp4_h_r_40_11904;
  wire seg_5_5_sp4_r_v_b_13_23157;
  wire seg_5_5_sp4_r_v_b_23_23167;
  wire seg_5_5_sp4_v_b_6_19209;
  wire seg_5_5_sp4_v_t_47_19705;
  wire seg_5_6_glb_netwk_0_5;
  wire seg_5_6_glb_netwk_7_12;
  wire seg_5_6_local_g0_0_23419;
  wire seg_5_6_local_g0_2_23421;
  wire seg_5_6_local_g0_3_23422;
  wire seg_5_6_local_g0_4_23423;
  wire seg_5_6_local_g0_5_23424;
  wire seg_5_6_local_g0_6_23425;
  wire seg_5_6_local_g0_7_23426;
  wire seg_5_6_local_g1_0_23427;
  wire seg_5_6_local_g2_1_23436;
  wire seg_5_6_local_g3_0_23443;
  wire seg_5_6_local_g3_2_23445;
  wire seg_5_6_local_g3_3_23446;
  wire seg_5_6_local_g3_5_23448;
  wire seg_5_6_lutff_1_out_19548;
  wire seg_5_6_lutff_2_out_19549;
  wire seg_5_6_lutff_3_out_19550;
  wire seg_5_6_lutff_4_out_19551;
  wire seg_5_6_lutff_5_out_19552;
  wire seg_5_6_lutff_6_out_19553;
  wire seg_5_6_neigh_op_bnl_0_15593;
  wire seg_5_6_sp12_h_r_11_1346;
  wire seg_5_6_sp4_h_l_37_7608;
  wire seg_5_6_sp4_h_l_41_7614;
  wire seg_5_6_sp4_h_r_10_23515;
  wire seg_5_6_sp4_h_r_2_23517;
  wire seg_5_6_sp4_h_r_30_15859;
  wire seg_5_6_sp4_h_r_33_15862;
  wire seg_5_6_sp4_r_v_b_19_23286;
  wire seg_5_6_sp4_r_v_b_21_23288;
  wire seg_5_6_sp4_v_b_0_19326;
  wire seg_5_6_sp4_v_b_10_19336;
  wire seg_5_6_sp4_v_b_12_19448;
  wire seg_5_6_sp4_v_b_13_19449;
  wire seg_5_6_sp4_v_b_14_19450;
  wire seg_5_6_sp4_v_b_15_19451;
  wire seg_5_6_sp4_v_b_26_19574;
  wire seg_5_6_sp4_v_b_8_19334;
  wire seg_5_6_sp4_v_t_38_19819;
  wire seg_5_6_sp4_v_t_40_19821;
  wire seg_5_6_sp4_v_t_42_19823;
  wire seg_5_6_sp4_v_t_47_19828;
  wire seg_5_7_glb_netwk_0_5;
  wire seg_5_7_glb_netwk_5_10;
  wire seg_5_7_local_g0_5_23547;
  wire seg_5_7_local_g0_6_23548;
  wire seg_5_7_local_g1_1_23551;
  wire seg_5_7_local_g1_3_23553;
  wire seg_5_7_local_g1_4_23554;
  wire seg_5_7_local_g1_5_23555;
  wire seg_5_7_local_g1_6_23556;
  wire seg_5_7_local_g3_1_23567;
  wire seg_5_7_local_g3_5_23571;
  wire seg_5_7_lutff_3_out_19673;
  wire seg_5_7_neigh_op_lft_1_15840;
  wire seg_5_7_neigh_op_lft_5_15844;
  wire seg_5_7_neigh_op_top_3_19796;
  wire seg_5_7_sp12_v_b_20_23389;
  wire seg_5_7_sp12_v_t_23_23635;
  wire seg_5_7_sp4_h_l_37_7755;
  wire seg_5_7_sp4_h_l_45_7765;
  wire seg_5_7_sp4_h_r_0_23636;
  wire seg_5_7_sp4_h_r_11_23639;
  wire seg_5_7_sp4_h_r_18_19814;
  wire seg_5_7_sp4_h_r_29_15981;
  wire seg_5_7_sp4_h_r_2_23640;
  wire seg_5_7_sp4_h_r_6_23644;
  wire seg_5_7_sp4_r_v_b_11_23289;
  wire seg_5_7_sp4_v_b_13_19572;
  wire seg_5_7_sp4_v_b_41_19822;
  wire seg_5_7_sp4_v_b_4_19453;
  wire seg_5_7_sp4_v_t_41_19945;
  wire seg_5_7_sp4_v_t_45_19949;
  wire seg_5_8_glb_netwk_0_5;
  wire seg_5_8_glb_netwk_4_9;
  wire seg_5_8_local_g0_3_23668;
  wire seg_5_8_local_g0_5_23670;
  wire seg_5_8_local_g0_6_23671;
  wire seg_5_8_local_g0_7_23672;
  wire seg_5_8_local_g1_1_23674;
  wire seg_5_8_local_g1_3_23676;
  wire seg_5_8_local_g1_5_23678;
  wire seg_5_8_local_g2_1_23682;
  wire seg_5_8_local_g2_3_23684;
  wire seg_5_8_local_g2_6_23687;
  wire seg_5_8_lutff_3_out_19796;
  wire seg_5_8_lutff_5_out_19798;
  wire seg_5_8_lutff_6_out_19799;
  wire seg_5_8_neigh_op_bnl_3_15842;
  wire seg_5_8_neigh_op_bot_3_19673;
  wire seg_5_8_sp12_v_b_23_23635;
  wire seg_5_8_sp4_h_l_39_7906;
  wire seg_5_8_sp4_h_l_41_7908;
  wire seg_5_8_sp4_h_l_43_7910;
  wire seg_5_8_sp4_h_l_44_7913;
  wire seg_5_8_sp4_h_l_47_7904;
  wire seg_5_8_sp4_h_r_11_23762;
  wire seg_5_8_sp4_h_r_14_19933;
  wire seg_5_8_sp4_h_r_1_23760;
  wire seg_5_8_sp4_h_r_20_19939;
  wire seg_5_8_sp4_h_r_3_23764;
  wire seg_5_8_sp4_h_r_5_23766;
  wire seg_5_8_sp4_h_r_6_23767;
  wire seg_5_8_sp4_h_r_7_23768;
  wire seg_5_8_sp4_h_r_8_23769;
  wire seg_5_8_sp4_h_r_9_23770;
  wire seg_5_8_sp4_r_v_b_1_23402;
  wire seg_5_8_sp4_r_v_b_23_23536;
  wire seg_5_8_sp4_v_b_15_19697;
  wire seg_5_8_sp4_v_b_22_19704;
  wire seg_5_8_sp4_v_b_2_19574;
  wire seg_5_8_sp4_v_b_33_19825;
  wire seg_5_8_sp4_v_t_37_20064;
  wire seg_5_8_sp4_v_t_39_20066;
  wire seg_5_8_sp4_v_t_43_20070;
  wire seg_5_8_sp4_v_t_46_20073;
  wire seg_5_8_sp4_v_t_47_20074;
  wire seg_5_9_glb_netwk_0_5;
  wire seg_5_9_glb_netwk_4_9;
  wire seg_5_9_local_g2_0_23804;
  wire seg_5_9_local_g2_1_23805;
  wire seg_5_9_local_g2_2_23806;
  wire seg_5_9_local_g2_3_23807;
  wire seg_5_9_local_g2_7_23811;
  wire seg_5_9_local_g3_0_23812;
  wire seg_5_9_local_g3_2_23814;
  wire seg_5_9_local_g3_5_23817;
  wire seg_5_9_neigh_op_rgt_0_23747;
  wire seg_5_9_neigh_op_rgt_2_23749;
  wire seg_5_9_neigh_op_rgt_5_23752;
  wire seg_5_9_neigh_op_tnr_0_23870;
  wire seg_5_9_neigh_op_tnr_1_23871;
  wire seg_5_9_neigh_op_tnr_2_23872;
  wire seg_5_9_neigh_op_tnr_3_23873;
  wire seg_5_9_neigh_op_tnr_7_23877;
  wire seg_5_9_sp12_h_r_10_1991;
  wire seg_5_9_sp4_h_l_36_8050;
  wire seg_5_9_sp4_h_l_46_8052;
  wire seg_5_9_sp4_h_r_0_23882;
  wire seg_5_9_sp4_h_r_16_20058;
  wire seg_5_9_sp4_h_r_20_20062;
  wire seg_5_9_sp4_h_r_22_20054;
  wire seg_5_9_sp4_r_v_b_25_23771;
  wire seg_5_9_sp4_r_v_b_27_23773;
  wire seg_5_9_sp4_r_v_b_29_23775;
  wire seg_5_9_sp4_r_v_b_33_23779;
  wire seg_5_9_sp4_r_v_b_35_23781;
  wire seg_5_9_sp4_v_b_0_19695;
  wire seg_5_9_sp4_v_b_36_20063;
  wire seg_5_9_sp4_v_b_38_20065;
  wire seg_5_9_sp4_v_b_40_20067;
  wire seg_5_9_sp4_v_b_42_20069;
  wire seg_5_9_sp4_v_b_44_20071;
  wire seg_5_9_sp4_v_b_46_20073;
  wire seg_5_9_sp4_v_b_4_19699;
  wire seg_5_9_sp4_v_b_9_19702;
  wire seg_5_9_sp4_v_t_37_20187;
  wire seg_5_9_sp4_v_t_39_20189;
  wire seg_5_9_sp4_v_t_41_20191;
  wire seg_5_9_sp4_v_t_46_20196;
  wire seg_6_0_span4_horz_r_6_22756;
  wire seg_6_0_span4_horz_r_8_18923;
  wire seg_6_0_span4_vert_0_22874;
  wire seg_6_0_span4_vert_28_22895;
  wire seg_6_10_glb_netwk_0_5;
  wire seg_6_10_local_g2_2_27569;
  wire seg_6_10_ram_RDATA_0_23877;
  wire seg_6_10_ram_RDATA_4_23873;
  wire seg_6_10_ram_RDATA_5_23872;
  wire seg_6_10_ram_RDATA_6_23871;
  wire seg_6_10_ram_RDATA_7_23870;
  wire seg_6_10_sp12_v_b_19_27318;
  wire seg_6_10_sp4_h_r_10_27627;
  wire seg_6_10_sp4_h_r_12_24006;
  wire seg_6_10_sp4_h_r_42_16352;
  wire seg_6_10_sp4_h_r_8_27635;
  wire seg_6_10_sp4_v_b_1_23648;
  wire seg_6_10_sp4_v_t_41_24145;
  wire seg_6_10_sp4_v_t_42_24146;
  wire seg_6_10_sp4_v_t_43_24147;
  wire seg_6_10_sp4_v_t_44_24148;
  wire seg_6_10_sp4_v_t_45_24149;
  wire seg_6_11_glb_netwk_0_5;
  wire seg_6_11_local_g0_2_27655;
  wire seg_6_11_local_g0_4_27657;
  wire seg_6_11_local_g0_6_27659;
  wire seg_6_11_local_g1_4_27665;
  wire seg_6_11_ram_RDATA_10_23998;
  wire seg_6_11_ram_RDATA_11_23997;
  wire seg_6_11_ram_RDATA_13_23995;
  wire seg_6_11_ram_RDATA_15_23993;
  wire seg_6_11_sp4_h_r_2_27731;
  wire seg_6_11_sp4_h_r_38_16471;
  wire seg_6_11_sp4_h_r_44_16477;
  wire seg_6_11_sp4_h_r_46_16469;
  wire seg_6_11_sp4_h_r_4_27733;
  wire seg_6_11_sp4_h_r_9_27738;
  wire seg_6_11_sp4_v_b_11_23781;
  wire seg_6_11_sp4_v_b_14_23896;
  wire seg_6_11_sp4_v_b_18_23900;
  wire seg_6_11_sp4_v_b_1_23771;
  wire seg_6_11_sp4_v_b_20_23902;
  wire seg_6_11_sp4_v_b_2_23774;
  wire seg_6_11_sp4_v_b_3_23773;
  wire seg_6_11_sp4_v_b_5_23775;
  wire seg_6_11_sp4_v_b_6_23778;
  wire seg_6_11_sp4_v_b_7_23777;
  wire seg_6_11_sp4_v_b_9_23779;
  wire seg_6_11_sp4_v_t_36_24263;
  wire seg_6_11_sp4_v_t_38_24265;
  wire seg_6_11_sp4_v_t_41_24268;
  wire seg_6_12_glb_netwk_0_5;
  wire seg_6_12_local_g1_3_27766;
  wire seg_6_12_ram_RDATA_3_24120;
  wire seg_6_12_ram_RDATA_7_24116;
  wire seg_6_12_sp4_h_r_0_27829;
  wire seg_6_12_sp4_h_r_11_27832;
  wire seg_6_12_sp4_h_r_14_24256;
  wire seg_6_12_sp4_h_r_28_20426;
  wire seg_6_12_sp4_h_r_34_20422;
  wire seg_6_12_sp4_h_r_6_27837;
  wire seg_6_12_sp4_v_b_10_23905;
  wire seg_6_12_sp4_v_b_1_23894;
  wire seg_6_12_sp4_v_b_2_23897;
  wire seg_6_12_sp4_v_b_36_24263;
  wire seg_6_12_sp4_v_b_38_24265;
  wire seg_6_12_sp4_v_b_6_23901;
  wire seg_6_12_sp4_v_t_42_24392;
  wire seg_6_12_sp4_v_t_45_24395;
  wire seg_6_13_sp4_h_l_36_12882;
  wire seg_6_13_sp4_h_l_47_12883;
  wire seg_6_13_sp4_v_b_2_24020;
  wire seg_6_13_sp4_v_b_4_24022;
  wire seg_6_13_sp4_v_b_7_24023;
  wire seg_6_13_sp4_v_t_39_24512;
  wire seg_6_14_sp4_v_b_1_24140;
  wire seg_6_14_sp4_v_t_37_24633;
  wire seg_6_14_sp4_v_t_43_24639;
  wire seg_6_15_sp4_v_b_10_24274;
  wire seg_6_15_sp4_v_b_2_24266;
  wire seg_6_15_sp4_v_b_5_24267;
  wire seg_6_16_sp4_v_t_40_24882;
  wire seg_6_18_sp4_v_t_37_25125;
  wire seg_6_19_sp12_v_t_23_28542;
  wire seg_6_1_sp4_h_l_36_11370;
  wire seg_6_1_sp4_h_l_38_11374;
  wire seg_6_1_sp4_h_l_42_11378;
  wire seg_6_1_sp4_h_l_44_11380;
  wire seg_6_1_sp4_h_r_9_26682;
  wire seg_6_1_sp4_v_b_0_22874;
  wire seg_6_20_sp4_v_t_40_25374;
  wire seg_6_22_sp4_v_t_41_25621;
  wire seg_6_24_sp4_v_t_40_25866;
  wire seg_6_25_sp4_h_r_1_29156;
  wire seg_6_26_sp4_v_t_36_26108;
  wire seg_6_28_sp4_v_t_40_26358;
  wire seg_6_29_sp4_h_r_3_29568;
  wire seg_6_2_sp4_h_l_37_11528;
  wire seg_6_2_sp4_h_l_43_11536;
  wire seg_6_2_sp4_h_l_45_11538;
  wire seg_6_2_sp4_v_t_45_23165;
  wire seg_6_30_sp4_v_t_40_29689;
  wire seg_6_31_local_g0_1_29708;
  wire seg_6_31_local_g0_1_29708_i1;
  wire seg_6_31_local_g0_1_29708_i2;
  wire seg_6_31_local_g0_1_29708_i3;
  wire seg_6_31_span12_vert_0_28542;
  wire seg_6_31_span4_vert_16_26358;
  wire seg_6_31_span4_vert_33_26481;
  wire seg_6_31_span4_vert_40_29689;
  wire seg_6_3_glb_netwk_0_5;
  wire seg_6_3_local_g0_2_26839;
  wire seg_6_3_local_g0_4_26841;
  wire seg_6_3_local_g0_6_26843;
  wire seg_6_3_local_g0_7_26844;
  wire seg_6_3_local_g1_2_26847;
  wire seg_6_3_local_g1_4_26849;
  wire seg_6_3_local_g1_5_26850;
  wire seg_6_3_local_g2_0_26853;
  wire seg_6_3_local_g2_2_26855;
  wire seg_6_3_local_g2_3_26856;
  wire seg_6_3_local_g2_7_26860;
  wire seg_6_3_local_g3_0_26861;
  wire seg_6_3_local_g3_1_26862;
  wire seg_6_3_local_g3_5_26866;
  wire seg_6_3_local_g3_6_26867;
  wire seg_6_3_neigh_op_lft_2_19180;
  wire seg_6_3_ram_RDATA_10_23014;
  wire seg_6_3_ram_RDATA_11_23013;
  wire seg_6_3_ram_RDATA_8_23016;
  wire seg_6_3_ram_RDATA_9_23015;
  wire seg_6_3_sp4_h_l_38_11656;
  wire seg_6_3_sp4_h_r_12_23145;
  wire seg_6_3_sp4_h_r_14_23149;
  wire seg_6_3_sp4_h_r_21_23154;
  wire seg_6_3_sp4_h_r_24_19313;
  wire seg_6_3_sp4_h_r_26_19317;
  wire seg_6_3_sp4_h_r_30_19321;
  wire seg_6_3_sp4_h_r_41_15488;
  wire seg_6_3_sp4_h_r_43_15490;
  wire seg_6_3_sp4_h_r_47_15484;
  wire seg_6_3_sp4_r_v_b_16_26718;
  wire seg_6_3_sp4_r_v_b_21_26723;
  wire seg_6_3_sp4_v_b_12_22904;
  wire seg_6_3_sp4_v_b_23_22916;
  wire seg_6_3_sp4_v_b_4_22895;
  wire seg_6_3_sp4_v_b_6_22898;
  wire seg_6_3_sp4_v_t_41_23284;
  wire seg_6_4_glb_netwk_0_5;
  wire seg_6_4_local_g0_0_26939;
  wire seg_6_4_local_g0_4_26943;
  wire seg_6_4_local_g0_5_26944;
  wire seg_6_4_local_g0_6_26945;
  wire seg_6_4_local_g1_2_26949;
  wire seg_6_4_local_g1_3_26950;
  wire seg_6_4_local_g1_4_26951;
  wire seg_6_4_local_g1_5_26952;
  wire seg_6_4_local_g2_0_26955;
  wire seg_6_4_local_g2_1_26956;
  wire seg_6_4_local_g2_2_26957;
  wire seg_6_4_local_g2_5_26960;
  wire seg_6_4_local_g2_6_26961;
  wire seg_6_4_local_g2_7_26962;
  wire seg_6_4_local_g3_1_26964;
  wire seg_6_4_local_g3_2_26965;
  wire seg_6_4_local_g3_5_26968;
  wire seg_6_4_local_g3_6_26969;
  wire seg_6_4_neigh_op_bnl_2_19180;
  wire seg_6_4_ram_RDATA_6_23133;
  wire seg_6_4_ram_RDATA_7_23132;
  wire seg_6_4_sp4_h_l_36_11775;
  wire seg_6_4_sp4_h_l_39_11778;
  wire seg_6_4_sp4_h_l_45_11784;
  wire seg_6_4_sp4_h_l_47_11776;
  wire seg_6_4_sp4_h_r_25_19437;
  wire seg_6_4_sp4_h_r_36_15606;
  wire seg_6_4_sp4_h_r_3_27018;
  wire seg_6_4_sp4_h_r_45_15615;
  wire seg_6_4_sp4_h_r_46_15608;
  wire seg_6_4_sp4_h_r_47_15607;
  wire seg_6_4_sp4_h_r_6_27021;
  wire seg_6_4_sp4_h_r_8_27023;
  wire seg_6_4_sp4_r_v_b_22_26831;
  wire seg_6_4_sp4_r_v_b_28_26928;
  wire seg_6_4_sp4_r_v_b_29_26927;
  wire seg_6_4_sp4_r_v_b_32_26932;
  wire seg_6_4_sp4_r_v_b_39_27028;
  wire seg_6_4_sp4_r_v_b_43_27032;
  wire seg_6_4_sp4_r_v_b_5_26718;
  wire seg_6_4_sp4_v_b_14_23035;
  wire seg_6_4_sp4_v_b_18_23039;
  wire seg_6_4_sp4_v_b_19_23040;
  wire seg_6_4_sp4_v_b_20_23041;
  wire seg_6_4_sp4_v_b_25_23156;
  wire seg_6_4_sp4_v_b_29_23160;
  wire seg_6_4_sp4_v_b_38_23281;
  wire seg_6_4_sp4_v_b_40_23283;
  wire seg_6_4_sp4_v_b_44_23287;
  wire seg_6_4_sp4_v_t_36_23402;
  wire seg_6_4_sp4_v_t_46_23412;
  wire seg_6_5_sp4_h_l_41_11903;
  wire seg_6_5_sp4_v_t_36_23525;
  wire seg_6_5_sp4_v_t_47_23536;
  wire seg_6_6_sp4_h_l_36_12021;
  wire seg_6_6_sp4_h_l_47_12022;
  wire seg_6_6_sp4_v_b_0_23157;
  wire seg_6_6_sp4_v_t_38_23650;
  wire seg_6_6_sp4_v_t_39_23651;
  wire seg_6_6_sp4_v_t_45_23657;
  wire seg_6_7_sp4_v_b_11_23289;
  wire seg_6_7_sp4_v_b_5_23283;
  wire seg_6_7_sp4_v_b_9_23287;
  wire seg_6_7_sp4_v_t_45_23780;
  wire seg_6_8_sp4_h_l_43_12274;
  wire seg_6_8_sp4_h_l_44_12277;
  wire seg_6_8_sp4_h_l_45_12276;
  wire seg_6_8_sp4_h_r_0_27421;
  wire seg_6_8_sp4_h_r_10_27423;
  wire seg_6_8_sp4_h_r_1_27422;
  wire seg_6_8_sp4_h_r_4_27427;
  wire seg_6_8_sp4_h_r_9_27432;
  wire seg_6_8_sp4_v_b_9_23410;
  wire seg_6_8_sp4_v_t_45_23903;
  wire seg_6_9_glb_netwk_0_5;
  wire seg_6_9_local_g2_2_27467;
  wire seg_6_9_local_g2_4_27469;
  wire seg_6_9_local_g2_6_27471;
  wire seg_6_9_local_g3_4_27477;
  wire seg_6_9_ram_RDATA_10_23752;
  wire seg_6_9_ram_RDATA_13_23749;
  wire seg_6_9_ram_RDATA_15_23747;
  wire seg_6_9_sp12_h_r_14_2002;
  wire seg_6_9_sp12_h_r_20_2012;
  wire seg_6_9_sp12_h_r_22_1992;
  wire seg_6_9_sp4_h_r_1_27524;
  wire seg_6_9_sp4_h_r_40_16227;
  wire seg_6_9_sp4_r_v_b_12_27331;
  wire seg_6_9_sp4_v_b_28_23776;
  wire seg_6_9_sp4_v_b_34_23782;
  wire seg_6_9_sp4_v_b_38_23896;
  wire seg_6_9_sp4_v_b_42_23900;
  wire seg_6_9_sp4_v_b_4_23530;
  wire seg_6_9_sp4_v_t_40_24021;
  wire seg_6_9_sp4_v_t_43_24024;
  wire seg_7_0_local_g1_7_29752;
  wire seg_7_0_span4_vert_15_26690;
  wire seg_7_10_glb_netwk_0_5;
  wire seg_7_10_glb_netwk_4_9;
  wire seg_7_10_local_g0_4_30946;
  wire seg_7_10_local_g1_0_30950;
  wire seg_7_10_local_g2_0_30958;
  wire seg_7_10_local_g2_1_30959;
  wire seg_7_10_local_g2_5_30963;
  wire seg_7_10_local_g3_1_30967;
  wire seg_7_10_local_g3_3_30969;
  wire seg_7_10_lutff_0_out_27481;
  wire seg_7_10_lutff_1_out_27482;
  wire seg_7_10_lutff_2_out_27483;
  wire seg_7_10_lutff_4_out_27485;
  wire seg_7_10_lutff_6_out_27487;
  wire seg_7_10_sp4_h_l_41_16349;
  wire seg_7_10_sp4_h_l_43_16351;
  wire seg_7_10_sp4_h_l_47_16345;
  wire seg_7_10_sp4_h_r_4_31042;
  wire seg_7_10_sp4_h_r_8_31046;
  wire seg_7_10_sp4_r_v_b_19_30809;
  wire seg_7_10_sp4_r_v_b_8_30688;
  wire seg_7_10_sp4_v_b_12_27433;
  wire seg_7_10_sp4_v_b_29_27539;
  wire seg_7_10_sp4_v_b_33_27543;
  wire seg_7_10_sp4_v_b_46_27647;
  wire seg_7_10_sp4_v_b_6_27338;
  wire seg_7_10_sp4_v_t_36_27739;
  wire seg_7_10_sp4_v_t_43_27746;
  wire seg_7_11_glb_netwk_0_5;
  wire seg_7_11_glb_netwk_4_9;
  wire seg_7_11_local_g0_6_31071;
  wire seg_7_11_local_g1_3_31076;
  wire seg_7_11_local_g1_6_31079;
  wire seg_7_11_local_g2_3_31084;
  wire seg_7_11_local_g2_5_31086;
  wire seg_7_11_local_g2_6_31087;
  wire seg_7_11_local_g3_2_31091;
  wire seg_7_11_local_g3_6_31095;
  wire seg_7_11_lutff_0_out_27583;
  wire seg_7_11_lutff_1_out_27584;
  wire seg_7_11_lutff_2_out_27585;
  wire seg_7_11_lutff_3_out_27586;
  wire seg_7_11_lutff_6_out_27589;
  wire seg_7_11_lutff_7_out_27590;
  wire seg_7_11_neigh_op_bot_6_27487;
  wire seg_7_11_sp4_h_l_36_16467;
  wire seg_7_11_sp4_h_r_30_24136;
  wire seg_7_11_sp4_h_r_37_20297;
  wire seg_7_11_sp4_h_r_42_20306;
  wire seg_7_11_sp4_h_r_46_20300;
  wire seg_7_11_sp4_h_r_4_31165;
  wire seg_7_11_sp4_h_r_8_31169;
  wire seg_7_11_sp4_r_v_b_11_30812;
  wire seg_7_11_sp4_v_b_10_27444;
  wire seg_7_11_sp4_v_b_26_27640;
  wire seg_7_11_sp4_v_b_3_27435;
  wire seg_7_11_sp4_v_b_40_27743;
  wire seg_7_11_sp4_v_b_7_27439;
  wire seg_7_11_sp4_v_t_39_27844;
  wire seg_7_11_sp4_v_t_45_27850;
  wire seg_7_12_local_g0_1_31189;
  wire seg_7_12_local_g0_2_31190;
  wire seg_7_12_local_g0_3_31191;
  wire seg_7_12_local_g0_4_31192;
  wire seg_7_12_local_g0_7_31195;
  wire seg_7_12_local_g1_0_31196;
  wire seg_7_12_local_g1_1_31197;
  wire seg_7_12_local_g1_2_31198;
  wire seg_7_12_local_g1_3_31199;
  wire seg_7_12_local_g1_5_31201;
  wire seg_7_12_local_g1_7_31203;
  wire seg_7_12_local_g2_3_31207;
  wire seg_7_12_local_g3_2_31214;
  wire seg_7_12_local_g3_5_31217;
  wire seg_7_12_lutff_1_out_27686;
  wire seg_7_12_lutff_2_out_27687;
  wire seg_7_12_lutff_3_out_27688;
  wire seg_7_12_lutff_4_out_27689;
  wire seg_7_12_lutff_5_out_27690;
  wire seg_7_12_lutff_6_out_27691;
  wire seg_7_12_lutff_7_out_27692;
  wire seg_7_12_neigh_op_bnr_1_31025;
  wire seg_7_12_neigh_op_bnr_3_31027;
  wire seg_7_12_neigh_op_bot_0_27583;
  wire seg_7_12_neigh_op_bot_1_27584;
  wire seg_7_12_neigh_op_bot_2_27585;
  wire seg_7_12_neigh_op_bot_3_27586;
  wire seg_7_12_neigh_op_bot_7_27590;
  wire seg_7_12_neigh_op_tnr_3_31273;
  wire seg_7_12_neigh_op_tnr_5_31275;
  wire seg_7_12_neigh_op_top_2_27789;
  wire seg_7_12_neigh_op_top_4_27791;
  wire seg_7_12_neigh_op_top_5_27792;
  wire seg_7_12_neigh_op_top_7_27794;
  wire seg_7_12_sp4_h_l_40_16596;
  wire seg_7_12_sp4_h_l_42_16598;
  wire seg_7_12_sp4_h_l_44_16600;
  wire seg_7_12_sp4_h_l_45_16599;
  wire seg_7_12_sp4_r_v_b_18_31054;
  wire seg_7_12_sp4_v_b_0_27536;
  wire seg_7_12_sp4_v_b_10_27546;
  wire seg_7_12_sp4_v_b_1_27535;
  wire seg_7_12_sp4_v_b_3_27537;
  wire seg_7_12_sp4_v_t_36_27943;
  wire seg_7_13_glb_netwk_0_5;
  wire seg_7_13_glb_netwk_4_9;
  wire seg_7_13_local_g0_1_31312;
  wire seg_7_13_local_g0_2_31313;
  wire seg_7_13_local_g0_3_31314;
  wire seg_7_13_local_g0_4_31315;
  wire seg_7_13_local_g1_0_31319;
  wire seg_7_13_local_g1_3_31322;
  wire seg_7_13_local_g2_4_31331;
  wire seg_7_13_local_g3_5_31340;
  wire seg_7_13_lutff_0_out_27787;
  wire seg_7_13_lutff_1_out_27788;
  wire seg_7_13_lutff_2_out_27789;
  wire seg_7_13_lutff_4_out_27791;
  wire seg_7_13_lutff_5_out_27792;
  wire seg_7_13_lutff_7_out_27794;
  wire seg_7_13_sp4_h_l_38_16717;
  wire seg_7_13_sp4_h_r_11_31408;
  wire seg_7_13_sp4_r_v_b_12_31171;
  wire seg_7_13_sp4_r_v_b_13_31172;
  wire seg_7_13_sp4_r_v_b_21_31180;
  wire seg_7_13_sp4_r_v_b_7_31054;
  wire seg_7_13_sp4_v_b_11_27647;
  wire seg_7_13_sp4_v_b_12_27739;
  wire seg_7_13_sp4_v_b_16_27743;
  wire seg_7_13_sp4_v_b_20_27747;
  wire seg_7_13_sp4_v_b_2_27640;
  wire seg_7_13_sp4_v_b_7_27643;
  wire seg_7_14_glb_netwk_0_5;
  wire seg_7_14_glb_netwk_4_9;
  wire seg_7_14_local_g1_2_31444;
  wire seg_7_14_local_g1_3_31445;
  wire seg_7_14_local_g1_6_31448;
  wire seg_7_14_local_g3_1_31459;
  wire seg_7_14_lutff_6_out_27895;
  wire seg_7_14_lutff_7_out_27896;
  wire seg_7_14_neigh_op_top_2_27993;
  wire seg_7_14_sp4_h_l_44_16846;
  wire seg_7_14_sp4_h_r_19_28041;
  wire seg_7_14_sp4_h_r_22_28036;
  wire seg_7_14_sp4_h_r_25_24498;
  wire seg_7_14_sp4_r_v_b_7_31177;
  wire seg_7_14_sp4_r_v_b_9_31179;
  wire seg_7_14_sp4_v_b_6_27746;
  wire seg_7_15_glb_netwk_0_5;
  wire seg_7_15_glb_netwk_4_9;
  wire seg_7_15_local_g0_0_31557;
  wire seg_7_15_local_g0_1_31558;
  wire seg_7_15_local_g0_2_31559;
  wire seg_7_15_local_g0_4_31561;
  wire seg_7_15_local_g0_5_31562;
  wire seg_7_15_local_g0_6_31563;
  wire seg_7_15_local_g0_7_31564;
  wire seg_7_15_local_g1_0_31565;
  wire seg_7_15_local_g1_1_31566;
  wire seg_7_15_local_g1_2_31567;
  wire seg_7_15_local_g1_3_31568;
  wire seg_7_15_local_g1_4_31569;
  wire seg_7_15_local_g1_5_31570;
  wire seg_7_15_local_g1_6_31571;
  wire seg_7_15_local_g1_7_31572;
  wire seg_7_15_local_g2_0_31573;
  wire seg_7_15_local_g2_1_31574;
  wire seg_7_15_local_g2_2_31575;
  wire seg_7_15_local_g2_4_31577;
  wire seg_7_15_local_g2_5_31578;
  wire seg_7_15_local_g3_1_31582;
  wire seg_7_15_local_g3_2_31583;
  wire seg_7_15_local_g3_3_31584;
  wire seg_7_15_local_g3_4_31585;
  wire seg_7_15_local_g3_5_31586;
  wire seg_7_15_lutff_2_out_27993;
  wire seg_7_15_neigh_op_bnr_6_31399;
  wire seg_7_15_neigh_op_top_0_28093;
  wire seg_7_15_sp12_v_b_2_30296;
  wire seg_7_15_sp12_v_b_4_30420;
  wire seg_7_15_sp4_h_l_40_16965;
  wire seg_7_15_sp4_h_l_42_16967;
  wire seg_7_15_sp4_h_r_16_28142;
  wire seg_7_15_sp4_h_r_21_28145;
  wire seg_7_15_sp4_h_r_23_28137;
  wire seg_7_15_sp4_h_r_29_24627;
  wire seg_7_15_sp4_h_r_40_20796;
  wire seg_7_15_sp4_r_v_b_10_31305;
  wire seg_7_15_sp4_r_v_b_11_31304;
  wire seg_7_15_sp4_r_v_b_17_31422;
  wire seg_7_15_sp4_r_v_b_19_31424;
  wire seg_7_15_sp4_r_v_b_20_31425;
  wire seg_7_15_sp4_r_v_b_21_31426;
  wire seg_7_15_sp4_r_v_b_31_31546;
  wire seg_7_15_sp4_r_v_b_3_31296;
  wire seg_7_15_sp4_r_v_b_7_31300;
  wire seg_7_15_sp4_r_v_b_9_31302;
  wire seg_7_15_sp4_v_b_10_27852;
  wire seg_7_15_sp4_v_b_12_27943;
  wire seg_7_15_sp4_v_b_13_27944;
  wire seg_7_15_sp4_v_b_14_27945;
  wire seg_7_15_sp4_v_b_16_27947;
  wire seg_7_15_sp4_v_b_17_27948;
  wire seg_7_15_sp4_v_b_18_27949;
  wire seg_7_15_sp4_v_b_1_27841;
  wire seg_7_15_sp4_v_b_23_27954;
  wire seg_7_15_sp4_v_b_2_27844;
  wire seg_7_15_sp4_v_b_4_27846;
  wire seg_7_15_sp4_v_b_8_27850;
  wire seg_7_16_glb_netwk_0_5;
  wire seg_7_16_glb_netwk_4_9;
  wire seg_7_16_local_g2_0_31696;
  wire seg_7_16_local_g2_3_31699;
  wire seg_7_16_local_g2_5_31701;
  wire seg_7_16_local_g3_5_31709;
  wire seg_7_16_local_g3_7_31711;
  wire seg_7_16_lutff_0_out_28093;
  wire seg_7_16_lutff_2_out_28095;
  wire seg_7_16_lutff_3_out_28096;
  wire seg_7_16_lutff_4_out_28097;
  wire seg_7_16_lutff_7_out_28100;
  wire seg_7_16_sp4_h_r_24_24743;
  wire seg_7_16_sp4_h_r_37_20912;
  wire seg_7_16_sp4_v_b_37_28250;
  wire seg_7_16_sp4_v_b_43_28256;
  wire seg_7_16_sp4_v_b_47_28260;
  wire seg_7_16_sp4_v_b_5_27947;
  wire seg_7_17_glb_netwk_0_5;
  wire seg_7_17_glb_netwk_4_9;
  wire seg_7_17_local_g0_2_31805;
  wire seg_7_17_local_g0_3_31806;
  wire seg_7_17_local_g0_4_31807;
  wire seg_7_17_local_g0_5_31808;
  wire seg_7_17_local_g1_0_31811;
  wire seg_7_17_local_g1_1_31812;
  wire seg_7_17_local_g1_2_31813;
  wire seg_7_17_local_g1_3_31814;
  wire seg_7_17_local_g1_5_31816;
  wire seg_7_17_local_g1_6_31817;
  wire seg_7_17_local_g1_7_31818;
  wire seg_7_17_local_g2_5_31824;
  wire seg_7_17_local_g3_5_31832;
  wire seg_7_17_local_g3_6_31833;
  wire seg_7_17_neigh_op_bot_2_28095;
  wire seg_7_17_neigh_op_bot_3_28096;
  wire seg_7_17_neigh_op_bot_4_28097;
  wire seg_7_17_neigh_op_bot_7_28100;
  wire seg_7_17_neigh_op_top_0_28297;
  wire seg_7_17_neigh_op_top_2_28299;
  wire seg_7_17_neigh_op_top_3_28300;
  wire seg_7_17_neigh_op_top_5_28302;
  wire seg_7_17_neigh_op_top_6_28303;
  wire seg_7_17_sp4_h_l_36_17205;
  wire seg_7_17_sp4_h_r_37_21035;
  wire seg_7_17_sp4_h_r_45_21045;
  wire seg_7_17_sp4_h_r_46_21038;
  wire seg_7_17_sp4_h_r_9_31908;
  wire seg_7_17_sp4_r_v_b_22_31673;
  wire seg_7_17_sp4_v_b_13_28148;
  wire seg_7_18_glb_netwk_0_5;
  wire seg_7_18_glb_netwk_4_9;
  wire seg_7_18_local_g0_6_31932;
  wire seg_7_18_local_g1_0_31934;
  wire seg_7_18_local_g1_3_31937;
  wire seg_7_18_local_g1_5_31939;
  wire seg_7_18_local_g3_4_31954;
  wire seg_7_18_local_g3_6_31956;
  wire seg_7_18_lutff_0_out_28297;
  wire seg_7_18_lutff_2_out_28299;
  wire seg_7_18_lutff_3_out_28300;
  wire seg_7_18_lutff_4_out_28301;
  wire seg_7_18_lutff_5_out_28302;
  wire seg_7_18_lutff_6_out_28303;
  wire seg_7_18_neigh_op_top_0_28399;
  wire seg_7_18_neigh_op_top_3_28402;
  wire seg_7_18_neigh_op_top_5_28404;
  wire seg_7_18_neigh_op_top_6_28405;
  wire seg_7_18_sp4_h_l_37_17327;
  wire seg_7_18_sp4_r_v_b_22_31796;
  wire seg_7_19_glb_netwk_0_5;
  wire seg_7_19_glb_netwk_4_9;
  wire seg_7_19_local_g2_0_32065;
  wire seg_7_19_local_g2_5_32070;
  wire seg_7_19_local_g2_7_32072;
  wire seg_7_19_local_g3_1_32074;
  wire seg_7_19_lutff_0_out_28399;
  wire seg_7_19_lutff_3_out_28402;
  wire seg_7_19_lutff_5_out_28404;
  wire seg_7_19_lutff_6_out_28405;
  wire seg_7_19_sp4_h_l_37_17450;
  wire seg_7_19_sp4_h_r_24_25112;
  wire seg_7_19_sp4_h_r_29_25119;
  wire seg_7_19_sp4_h_r_33_25123;
  wire seg_7_19_sp4_r_v_b_15_31912;
  wire seg_7_1_glb_netwk_0_5;
  wire seg_7_1_glb_netwk_4_9;
  wire seg_7_1_local_g3_4_29823;
  wire seg_7_1_lutff_1_out_26554;
  wire seg_7_1_sp4_h_l_43_15208;
  wire seg_7_1_sp4_h_r_8_29903;
  wire seg_7_1_sp4_r_v_b_44_29944;
  wire seg_7_2_glb_netwk_0_5;
  wire seg_7_2_glb_netwk_4_9;
  wire seg_7_2_local_g0_3_29961;
  wire seg_7_2_local_g2_6_29980;
  wire seg_7_2_local_g3_1_29983;
  wire seg_7_2_lutff_2_out_26631;
  wire seg_7_2_lutff_3_out_26632;
  wire seg_7_2_lutff_4_out_26633;
  wire seg_7_2_sp4_h_l_41_15365;
  wire seg_7_2_sp4_h_l_45_15369;
  wire seg_7_2_sp4_h_r_4_30058;
  wire seg_7_2_sp4_h_r_7_30061;
  wire seg_7_2_sp4_h_r_9_30063;
  wire seg_7_2_sp4_v_b_25_26713;
  wire seg_7_2_sp4_v_b_30_26721;
  wire seg_7_3_glb_netwk_0_5;
  wire seg_7_3_glb_netwk_4_9;
  wire seg_7_3_local_g0_0_30081;
  wire seg_7_3_local_g1_2_30091;
  wire seg_7_3_local_g2_7_30104;
  wire seg_7_3_local_g3_7_30112;
  wire seg_7_3_lutff_2_out_26769;
  wire seg_7_3_neigh_op_top_0_26869;
  wire seg_7_3_sp4_h_r_0_30175;
  wire seg_7_3_sp4_h_r_22_26914;
  wire seg_7_3_sp4_h_r_3_30180;
  wire seg_7_3_sp4_h_r_5_30182;
  wire seg_7_3_sp4_h_r_6_30183;
  wire seg_7_3_sp4_h_r_8_30185;
  wire seg_7_3_sp4_h_r_9_30186;
  wire seg_7_3_sp4_r_v_b_15_29938;
  wire seg_7_3_sp4_r_v_b_23_29947;
  wire seg_7_4_glb_netwk_0_5;
  wire seg_7_4_glb_netwk_4_9;
  wire seg_7_4_local_g0_4_30208;
  wire seg_7_4_local_g0_7_30211;
  wire seg_7_4_local_g2_1_30221;
  wire seg_7_4_local_g2_4_30224;
  wire seg_7_4_local_g2_5_30225;
  wire seg_7_4_local_g3_4_30232;
  wire seg_7_4_local_g3_7_30235;
  wire seg_7_4_lutff_0_out_26869;
  wire seg_7_4_lutff_1_out_26870;
  wire seg_7_4_lutff_2_out_26871;
  wire seg_7_4_neigh_op_rgt_4_30167;
  wire seg_7_4_sp4_h_l_42_15614;
  wire seg_7_4_sp4_h_r_0_30298;
  wire seg_7_4_sp4_h_r_12_27014;
  wire seg_7_4_sp4_h_r_28_23273;
  wire seg_7_4_sp4_h_r_2_30302;
  wire seg_7_4_sp4_h_r_3_30303;
  wire seg_7_4_sp4_h_r_42_19445;
  wire seg_7_4_sp4_h_r_45_19446;
  wire seg_7_4_sp4_h_r_6_30306;
  wire seg_7_4_sp4_h_r_7_30307;
  wire seg_7_4_sp4_h_r_8_30308;
  wire seg_7_4_sp4_r_v_b_23_30075;
  wire seg_7_4_sp4_r_v_b_27_30189;
  wire seg_7_4_sp4_r_v_b_47_30321;
  wire seg_7_4_sp4_v_b_6_26721;
  wire seg_7_4_sp4_v_t_36_27127;
  wire seg_7_5_glb_netwk_0_5;
  wire seg_7_5_glb_netwk_3_8;
  wire seg_7_5_local_g0_2_30329;
  wire seg_7_5_local_g0_6_30333;
  wire seg_7_5_local_g1_1_30336;
  wire seg_7_5_local_g1_2_30337;
  wire seg_7_5_local_g1_6_30341;
  wire seg_7_5_local_g1_7_30342;
  wire seg_7_5_local_g2_0_30343;
  wire seg_7_5_local_g2_3_30346;
  wire seg_7_5_local_g2_5_30348;
  wire seg_7_5_local_g2_7_30350;
  wire seg_7_5_local_g3_3_30354;
  wire seg_7_5_local_g3_4_30355;
  wire seg_7_5_local_g3_7_30358;
  wire seg_7_5_lutff_1_out_26972;
  wire seg_7_5_lutff_2_out_26973;
  wire seg_7_5_lutff_3_out_26974;
  wire seg_7_5_lutff_5_out_26976;
  wire seg_7_5_lutff_7_out_26978;
  wire seg_7_5_neigh_op_bot_2_26871;
  wire seg_7_5_neigh_op_rgt_3_30289;
  wire seg_7_5_neigh_op_rgt_7_30293;
  wire seg_7_5_sp4_h_l_36_15729;
  wire seg_7_5_sp4_h_l_42_15737;
  wire seg_7_5_sp4_h_l_44_15739;
  wire seg_7_5_sp4_h_l_46_15731;
  wire seg_7_5_sp4_h_r_10_30423;
  wire seg_7_5_sp4_h_r_14_27120;
  wire seg_7_5_sp4_h_r_22_27118;
  wire seg_7_5_sp4_h_r_24_23390;
  wire seg_7_5_sp4_h_r_47_19561;
  wire seg_7_5_sp4_h_r_9_30432;
  wire seg_7_5_sp4_r_v_b_19_30194;
  wire seg_7_5_sp4_r_v_b_25_30310;
  wire seg_7_5_sp4_v_b_24_27026;
  wire seg_7_5_sp4_v_b_28_27030;
  wire seg_7_5_sp4_v_b_44_27135;
  wire seg_7_5_sp4_v_b_45_27136;
  wire seg_7_6_glb_netwk_0_5;
  wire seg_7_6_glb_netwk_4_9;
  wire seg_7_6_local_g0_3_30453;
  wire seg_7_6_local_g0_5_30455;
  wire seg_7_6_local_g1_1_30459;
  wire seg_7_6_local_g1_2_30460;
  wire seg_7_6_local_g1_3_30461;
  wire seg_7_6_local_g1_5_30463;
  wire seg_7_6_local_g3_2_30476;
  wire seg_7_6_local_g3_3_30477;
  wire seg_7_6_local_g3_4_30478;
  wire seg_7_6_local_g3_7_30481;
  wire seg_7_6_lutff_2_out_27075;
  wire seg_7_6_lutff_3_out_27076;
  wire seg_7_6_lutff_7_out_27080;
  wire seg_7_6_neigh_op_bot_1_26972;
  wire seg_7_6_neigh_op_bot_2_26973;
  wire seg_7_6_neigh_op_bot_3_26974;
  wire seg_7_6_neigh_op_bot_5_26976;
  wire seg_7_6_sp4_h_l_40_15858;
  wire seg_7_6_sp4_h_l_43_15859;
  wire seg_7_6_sp4_h_l_45_15861;
  wire seg_7_6_sp4_h_r_13_27217;
  wire seg_7_6_sp4_h_r_26_23517;
  wire seg_7_6_sp4_h_r_27_23518;
  wire seg_7_6_sp4_h_r_34_23515;
  wire seg_7_6_sp4_h_r_40_19689;
  wire seg_7_6_sp4_h_r_44_19693;
  wire seg_7_6_sp4_v_b_12_27025;
  wire seg_7_6_sp4_v_b_42_27235;
  wire seg_7_6_sp4_v_b_44_27237;
  wire seg_7_7_glb_netwk_0_5;
  wire seg_7_7_glb_netwk_4_9;
  wire seg_7_7_local_g0_2_30575;
  wire seg_7_7_local_g0_3_30576;
  wire seg_7_7_local_g0_6_30579;
  wire seg_7_7_local_g0_7_30580;
  wire seg_7_7_local_g1_3_30584;
  wire seg_7_7_local_g2_2_30591;
  wire seg_7_7_local_g2_3_30592;
  wire seg_7_7_local_g3_4_30601;
  wire seg_7_7_local_g3_7_30604;
  wire seg_7_7_lutff_0_out_27175;
  wire seg_7_7_lutff_1_out_27176;
  wire seg_7_7_lutff_2_out_27177;
  wire seg_7_7_lutff_3_out_27178;
  wire seg_7_7_lutff_6_out_27181;
  wire seg_7_7_lutff_7_out_27182;
  wire seg_7_7_sp4_h_l_37_15974;
  wire seg_7_7_sp4_h_r_10_30669;
  wire seg_7_7_sp4_h_r_11_30670;
  wire seg_7_7_sp4_h_r_22_27322;
  wire seg_7_7_sp4_h_r_24_23636;
  wire seg_7_7_sp4_h_r_26_23640;
  wire seg_7_7_sp4_h_r_28_23642;
  wire seg_7_7_sp4_h_r_39_19809;
  wire seg_7_7_sp4_h_r_3_30672;
  wire seg_7_7_sp4_v_b_11_27035;
  wire seg_7_7_sp4_v_b_1_27025;
  wire seg_7_7_sp4_v_b_2_27028;
  wire seg_7_7_sp4_v_b_6_27032;
  wire seg_7_7_sp4_v_t_40_27437;
  wire seg_7_7_sp4_v_t_41_27438;
  wire seg_7_7_sp4_v_t_45_27442;
  wire seg_7_7_sp4_v_t_46_27443;
  wire seg_7_8_glb_netwk_0_5;
  wire seg_7_8_glb_netwk_4_9;
  wire seg_7_8_local_g0_0_30696;
  wire seg_7_8_local_g0_6_30702;
  wire seg_7_8_local_g1_0_30704;
  wire seg_7_8_local_g2_0_30712;
  wire seg_7_8_local_g2_6_30718;
  wire seg_7_8_local_g3_0_30720;
  wire seg_7_8_local_g3_4_30724;
  wire seg_7_8_local_g3_6_30726;
  wire seg_7_8_lutff_0_out_27277;
  wire seg_7_8_lutff_1_out_27278;
  wire seg_7_8_lutff_2_out_27279;
  wire seg_7_8_lutff_4_out_27281;
  wire seg_7_8_lutff_5_out_27282;
  wire seg_7_8_lutff_6_out_27283;
  wire seg_7_8_lutff_7_out_27284;
  wire seg_7_8_neigh_op_bot_0_27175;
  wire seg_7_8_neigh_op_bot_6_27181;
  wire seg_7_8_sp4_h_l_36_16098;
  wire seg_7_8_sp4_h_l_37_16097;
  wire seg_7_8_sp4_h_r_24_23759;
  wire seg_7_8_sp4_h_r_32_23769;
  wire seg_7_8_sp4_h_r_38_19933;
  wire seg_7_8_sp4_h_r_44_19939;
  wire seg_7_8_sp4_v_b_2_27130;
  wire seg_7_8_sp4_v_b_30_27338;
  wire seg_7_8_sp4_v_b_38_27435;
  wire seg_7_8_sp4_v_b_9_27135;
  wire seg_7_9_glb_netwk_0_5;
  wire seg_7_9_glb_netwk_5_10;
  wire seg_7_9_local_g0_1_30820;
  wire seg_7_9_local_g1_1_30828;
  wire seg_7_9_local_g1_3_30830;
  wire seg_7_9_local_g1_4_30831;
  wire seg_7_9_local_g2_1_30836;
  wire seg_7_9_local_g2_6_30841;
  wire seg_7_9_local_g3_5_30848;
  wire seg_7_9_sp12_v_b_14_30296;
  wire seg_7_9_sp12_v_b_16_30420;
  wire seg_7_9_sp4_h_r_12_27524;
  wire seg_7_9_sp4_h_r_17_27529;
  wire seg_7_9_sp4_h_r_19_27531;
  wire seg_7_9_sp4_h_r_24_23882;
  wire seg_7_9_sp4_h_r_25_23883;
  wire seg_7_9_sp4_r_v_b_38_30927;
  wire seg_7_9_sp4_v_b_17_27336;
  wire seg_7_9_sp4_v_b_20_27339;
  wire seg_7_9_sp4_v_b_34_27444;
  wire seg_7_9_sp4_v_b_36_27535;
  wire seg_7_9_sp4_v_b_38_27537;
  wire seg_7_9_sp4_v_b_45_27544;
  wire seg_7_9_sp4_v_b_7_27235;
  wire seg_8_0_local_g0_4_33572;
  wire seg_8_0_span4_vert_36_29935;
  wire seg_8_10_glb_netwk_0_5;
  wire seg_8_10_local_g0_0_34773;
  wire seg_8_10_local_g1_7_34788;
  wire seg_8_10_local_g2_2_34791;
  wire seg_8_10_sp4_h_l_41_20180;
  wire seg_8_10_sp4_h_l_43_20182;
  wire seg_8_10_sp4_h_r_23_31038;
  wire seg_8_10_sp4_h_r_4_34873;
  wire seg_8_10_sp4_h_r_8_34877;
  wire seg_8_10_sp4_v_b_1_30679;
  wire seg_8_10_sp4_v_b_26_30928;
  wire seg_8_10_sp4_v_b_34_30936;
  wire seg_8_10_sp4_v_b_36_31048;
  wire seg_8_10_sp4_v_b_3_30681;
  wire seg_8_10_sp4_v_b_5_30683;
  wire seg_8_10_sp4_v_t_37_31172;
  wire seg_8_10_sp4_v_t_42_31177;
  wire seg_8_11_glb_netwk_0_5;
  wire seg_8_11_glb_netwk_4_9;
  wire seg_8_11_local_g1_0_34904;
  wire seg_8_11_local_g1_2_34906;
  wire seg_8_11_local_g1_4_34908;
  wire seg_8_11_local_g2_4_34916;
  wire seg_8_11_local_g2_6_34918;
  wire seg_8_11_local_g3_0_34920;
  wire seg_8_11_local_g3_2_34922;
  wire seg_8_11_local_g3_6_34926;
  wire seg_8_11_lutff_0_out_31024;
  wire seg_8_11_lutff_1_out_31025;
  wire seg_8_11_lutff_2_out_31026;
  wire seg_8_11_lutff_3_out_31027;
  wire seg_8_11_lutff_4_out_31028;
  wire seg_8_11_lutff_6_out_31030;
  wire seg_8_11_sp12_v_b_0_33605;
  wire seg_8_11_sp4_h_l_43_20305;
  wire seg_8_11_sp4_h_l_44_20308;
  wire seg_8_11_sp4_h_l_45_20307;
  wire seg_8_11_sp4_h_r_0_34990;
  wire seg_8_11_sp4_h_r_14_31164;
  wire seg_8_11_sp4_h_r_1_34991;
  wire seg_8_11_sp4_h_r_38_24133;
  wire seg_8_11_sp4_h_r_4_34996;
  wire seg_8_11_sp4_h_r_5_34997;
  wire seg_8_11_sp4_h_r_6_34998;
  wire seg_8_11_sp4_r_v_b_15_34759;
  wire seg_8_11_sp4_v_b_0_30803;
  wire seg_8_11_sp4_v_b_10_30813;
  wire seg_8_11_sp4_v_b_14_30927;
  wire seg_8_11_sp4_v_b_1_30802;
  wire seg_8_11_sp4_v_b_26_31051;
  wire seg_8_11_sp4_v_b_2_30805;
  wire seg_8_11_sp4_v_b_44_31179;
  wire seg_8_11_sp4_v_b_9_30810;
  wire seg_8_11_sp4_v_t_42_31300;
  wire seg_8_11_sp4_v_t_46_31304;
  wire seg_8_12_glb_netwk_0_5;
  wire seg_8_12_glb_netwk_4_9;
  wire seg_8_12_local_g0_2_35021;
  wire seg_8_12_local_g0_4_35023;
  wire seg_8_12_local_g1_1_35028;
  wire seg_8_12_local_g1_3_35030;
  wire seg_8_12_local_g1_5_35032;
  wire seg_8_12_local_g1_6_35033;
  wire seg_8_12_local_g1_7_35034;
  wire seg_8_12_local_g2_0_35035;
  wire seg_8_12_local_g2_5_35040;
  wire seg_8_12_neigh_op_lft_1_27686;
  wire seg_8_12_neigh_op_lft_2_27687;
  wire seg_8_12_neigh_op_lft_3_27688;
  wire seg_8_12_neigh_op_lft_4_27689;
  wire seg_8_12_neigh_op_lft_5_27690;
  wire seg_8_12_neigh_op_lft_6_27691;
  wire seg_8_12_neigh_op_lft_7_27692;
  wire seg_8_12_neigh_op_rgt_5_34983;
  wire seg_8_12_neigh_op_tnl_0_27787;
  wire seg_8_12_sp12_v_b_19_34743;
  wire seg_8_12_sp4_h_l_42_20429;
  wire seg_8_12_sp4_h_l_46_20423;
  wire seg_8_12_sp4_h_r_10_35115;
  wire seg_8_12_sp4_h_r_2_35117;
  wire seg_8_12_sp4_h_r_5_35120;
  wire seg_8_12_sp4_h_r_6_35121;
  wire seg_8_12_sp4_h_r_7_35122;
  wire seg_8_12_sp4_h_r_8_35123;
  wire seg_8_12_sp4_h_r_9_35124;
  wire seg_8_12_sp4_r_v_b_15_34882;
  wire seg_8_12_sp4_v_b_10_30936;
  wire seg_8_12_sp4_v_b_4_30930;
  wire seg_8_12_sp4_v_b_5_30929;
  wire seg_8_12_sp4_v_b_6_30932;
  wire seg_8_12_sp4_v_b_9_30933;
  wire seg_8_13_glb_netwk_0_5;
  wire seg_8_13_glb_netwk_4_9;
  wire seg_8_13_local_g1_4_35154;
  wire seg_8_13_local_g2_0_35158;
  wire seg_8_13_local_g2_3_35161;
  wire seg_8_13_local_g3_2_35168;
  wire seg_8_13_local_g3_4_35170;
  wire seg_8_13_local_g3_6_35172;
  wire seg_8_13_local_g3_7_35173;
  wire seg_8_13_lutff_0_out_31270;
  wire seg_8_13_lutff_3_out_31273;
  wire seg_8_13_lutff_4_out_31274;
  wire seg_8_13_lutff_5_out_31275;
  wire seg_8_13_lutff_6_out_31276;
  wire seg_8_13_neigh_op_tnl_7_27896;
  wire seg_8_13_sp4_h_l_37_20543;
  wire seg_8_13_sp4_h_r_28_27937;
  wire seg_8_13_sp4_h_r_43_24382;
  wire seg_8_13_sp4_r_v_b_31_35131;
  wire seg_8_13_sp4_v_b_0_31049;
  wire seg_8_13_sp4_v_b_11_31058;
  wire seg_8_13_sp4_v_b_1_31048;
  wire seg_8_13_sp4_v_b_26_31297;
  wire seg_8_13_sp4_v_b_2_31051;
  wire seg_8_13_sp4_v_b_4_31053;
  wire seg_8_13_sp4_v_b_5_31052;
  wire seg_8_13_sp4_v_b_9_31056;
  wire seg_8_13_sp4_v_t_42_31546;
  wire seg_8_14_glb_netwk_0_5;
  wire seg_8_14_glb_netwk_3_8;
  wire seg_8_14_local_g0_4_35269;
  wire seg_8_14_local_g1_0_35273;
  wire seg_8_14_local_g1_3_35276;
  wire seg_8_14_local_g2_0_35281;
  wire seg_8_14_local_g2_1_35282;
  wire seg_8_14_lutff_0_out_31393;
  wire seg_8_14_lutff_6_out_31399;
  wire seg_8_14_sp4_h_r_6_35367;
  wire seg_8_14_sp4_h_r_7_35368;
  wire seg_8_14_sp4_r_v_b_27_35250;
  wire seg_8_14_sp4_r_v_b_9_35010;
  wire seg_8_14_sp4_v_b_12_31294;
  wire seg_8_14_sp4_v_b_16_31298;
  wire seg_8_14_sp4_v_b_6_31178;
  wire seg_8_15_glb_netwk_0_5;
  wire seg_8_15_local_g0_0_35388;
  wire seg_8_15_local_g0_2_35390;
  wire seg_8_15_local_g0_3_35391;
  wire seg_8_15_local_g0_4_35392;
  wire seg_8_15_local_g0_6_35394;
  wire seg_8_15_local_g1_0_35396;
  wire seg_8_15_local_g1_1_35397;
  wire seg_8_15_local_g1_3_35399;
  wire seg_8_15_local_g1_4_35400;
  wire seg_8_15_local_g1_5_35401;
  wire seg_8_15_local_g1_6_35402;
  wire seg_8_15_local_g1_7_35403;
  wire seg_8_15_local_g2_0_35404;
  wire seg_8_15_local_g2_1_35405;
  wire seg_8_15_local_g2_2_35406;
  wire seg_8_15_local_g2_3_35407;
  wire seg_8_15_local_g2_6_35410;
  wire seg_8_15_local_g3_1_35413;
  wire seg_8_15_local_g3_2_35414;
  wire seg_8_15_local_g3_3_35415;
  wire seg_8_15_local_g3_4_35416;
  wire seg_8_15_local_g3_5_35417;
  wire seg_8_15_local_g3_7_35419;
  wire seg_8_15_neigh_op_bnr_0_35224;
  wire seg_8_15_neigh_op_rgt_0_35347;
  wire seg_8_15_neigh_op_rgt_1_35348;
  wire seg_8_15_neigh_op_rgt_3_35350;
  wire seg_8_15_neigh_op_rgt_4_35351;
  wire seg_8_15_neigh_op_rgt_5_35352;
  wire seg_8_15_neigh_op_rgt_6_35353;
  wire seg_8_15_neigh_op_rgt_7_35354;
  wire seg_8_15_sp4_h_r_0_35482;
  wire seg_8_15_sp4_h_r_11_35485;
  wire seg_8_15_sp4_h_r_12_31652;
  wire seg_8_15_sp4_h_r_19_31659;
  wire seg_8_15_sp4_h_r_1_35483;
  wire seg_8_15_sp4_h_r_23_31653;
  wire seg_8_15_sp4_h_r_26_28139;
  wire seg_8_15_sp4_h_r_4_35488;
  wire seg_8_15_sp4_r_v_b_11_35135;
  wire seg_8_15_sp4_r_v_b_15_35251;
  wire seg_8_15_sp4_r_v_b_39_35497;
  wire seg_8_15_sp4_r_v_b_3_35127;
  wire seg_8_15_sp4_r_v_b_41_35499;
  wire seg_8_15_sp4_r_v_b_4_35130;
  wire seg_8_15_sp4_r_v_b_5_35129;
  wire seg_8_15_sp4_v_b_0_31295;
  wire seg_8_15_sp4_v_b_12_31417;
  wire seg_8_15_sp4_v_b_18_31423;
  wire seg_8_15_sp4_v_b_22_31427;
  wire seg_8_15_sp4_v_b_25_31540;
  wire seg_8_15_sp4_v_b_42_31669;
  wire seg_8_15_sp4_v_b_6_31301;
  wire seg_8_16_glb_netwk_0_5;
  wire seg_8_16_glb_netwk_4_9;
  wire seg_8_16_local_g0_2_35513;
  wire seg_8_16_local_g0_4_35515;
  wire seg_8_16_local_g1_0_35519;
  wire seg_8_16_local_g1_3_35522;
  wire seg_8_16_local_g1_5_35524;
  wire seg_8_16_local_g1_6_35525;
  wire seg_8_16_local_g1_7_35526;
  wire seg_8_16_local_g2_1_35528;
  wire seg_8_16_local_g2_3_35530;
  wire seg_8_16_local_g2_6_35533;
  wire seg_8_16_local_g3_0_35535;
  wire seg_8_16_local_g3_1_35536;
  wire seg_8_16_sp12_v_b_3_34251;
  wire seg_8_16_sp4_h_r_22_31777;
  wire seg_8_16_sp4_h_r_3_35610;
  wire seg_8_16_sp4_h_r_4_35611;
  wire seg_8_16_sp4_r_v_b_13_35372;
  wire seg_8_16_sp4_r_v_b_14_35373;
  wire seg_8_16_sp4_r_v_b_16_35375;
  wire seg_8_16_sp4_r_v_b_17_35376;
  wire seg_8_16_sp4_r_v_b_19_35378;
  wire seg_8_16_sp4_r_v_b_7_35254;
  wire seg_8_16_sp4_r_v_b_9_35256;
  wire seg_8_16_sp4_v_b_15_31543;
  wire seg_8_16_sp4_v_b_16_31544;
  wire seg_8_16_sp4_v_b_20_31548;
  wire seg_8_16_sp4_v_b_21_31549;
  wire seg_8_16_sp4_v_b_2_31420;
  wire seg_8_17_sp4_h_r_0_35728;
  wire seg_8_17_sp4_h_r_6_35736;
  wire seg_8_18_sp4_h_l_46_21161;
  wire seg_8_18_sp4_v_b_9_31671;
  wire seg_8_19_sp12_v_t_23_35973;
  wire seg_8_19_sp4_h_l_40_21288;
  wire seg_8_1_glb_netwk_0_5;
  wire seg_8_1_glb_netwk_4_9;
  wire seg_8_1_local_g1_1_33635;
  wire seg_8_1_local_g2_2_33644;
  wire seg_8_1_local_g2_4_33646;
  wire seg_8_1_local_g2_6_33648;
  wire seg_8_1_local_g3_2_33652;
  wire seg_8_1_lutff_2_out_29755;
  wire seg_8_1_lutff_3_out_29756;
  wire seg_8_1_lutff_5_out_29758;
  wire seg_8_1_lutff_6_out_29759;
  wire seg_8_1_lutff_7_out_29760;
  wire seg_8_1_neigh_op_lft_1_26554;
  wire seg_8_1_neigh_op_tnl_2_26631;
  wire seg_8_1_neigh_op_tnl_4_26633;
  wire seg_8_1_sp4_h_r_2_33728;
  wire seg_8_20_sp4_h_l_39_21408;
  wire seg_8_21_sp12_v_t_23_36219;
  wire seg_8_22_sp4_v_b_0_32156;
  wire seg_8_2_glb_netwk_0_5;
  wire seg_8_2_glb_netwk_4_9;
  wire seg_8_2_local_g2_7_33812;
  wire seg_8_2_local_g3_0_33813;
  wire seg_8_2_local_g3_5_33818;
  wire seg_8_2_lutff_0_out_29881;
  wire seg_8_2_sp4_h_r_4_33889;
  wire seg_8_2_sp4_r_v_b_29_33771;
  wire seg_8_2_sp4_v_b_29_29940;
  wire seg_8_2_sp4_v_b_39_30067;
  wire seg_8_2_sp4_v_t_37_30188;
  wire seg_8_31_span12_vert_0_35973;
  wire seg_8_31_span12_vert_4_36219;
  wire seg_8_3_glb_netwk_0_5;
  wire seg_8_3_local_g0_2_33914;
  wire seg_8_3_local_g0_5_33917;
  wire seg_8_3_local_g0_6_33918;
  wire seg_8_3_local_g2_3_33931;
  wire seg_8_3_local_g2_5_33933;
  wire seg_8_3_local_g2_6_33934;
  wire seg_8_3_local_g2_7_33935;
  wire seg_8_3_local_g3_1_33937;
  wire seg_8_3_local_g3_5_33941;
  wire seg_8_3_lutff_5_out_30045;
  wire seg_8_3_lutff_7_out_30047;
  wire seg_8_3_neigh_op_bnr_6_33718;
  wire seg_8_3_sp4_h_l_41_19319;
  wire seg_8_3_sp4_h_r_11_34009;
  wire seg_8_3_sp4_h_r_16_30182;
  wire seg_8_3_sp4_h_r_30_26919;
  wire seg_8_3_sp4_r_v_b_11_33765;
  wire seg_8_3_sp4_r_v_b_13_33767;
  wire seg_8_3_sp4_r_v_b_17_33772;
  wire seg_8_3_sp4_v_b_18_29942;
  wire seg_8_3_sp4_v_b_28_30069;
  wire seg_8_3_sp4_v_b_37_30188;
  wire seg_8_3_sp4_v_t_36_30310;
  wire seg_8_3_sp4_v_t_47_30321;
  wire seg_8_4_glb_netwk_0_5;
  wire seg_8_4_glb_netwk_4_9;
  wire seg_8_4_local_g0_3_34038;
  wire seg_8_4_local_g0_5_34040;
  wire seg_8_4_local_g1_2_34045;
  wire seg_8_4_local_g2_2_34053;
  wire seg_8_4_local_g2_4_34055;
  wire seg_8_4_local_g2_5_34056;
  wire seg_8_4_local_g3_5_34064;
  wire seg_8_4_lutff_2_out_30165;
  wire seg_8_4_lutff_4_out_30167;
  wire seg_8_4_lutff_5_out_30168;
  wire seg_8_4_sp4_h_l_38_19441;
  wire seg_8_4_sp4_h_l_39_19440;
  wire seg_8_4_sp4_h_l_40_19443;
  wire seg_8_4_sp4_h_l_41_19442;
  wire seg_8_4_sp4_h_l_44_19447;
  wire seg_8_4_sp4_h_r_11_34132;
  wire seg_8_4_sp4_h_r_16_30305;
  wire seg_8_4_sp4_h_r_1_34130;
  wire seg_8_4_sp4_h_r_22_30301;
  wire seg_8_4_sp4_h_r_29_27020;
  wire seg_8_4_sp4_h_r_2_34133;
  wire seg_8_4_sp4_h_r_37_23267;
  wire seg_8_4_sp4_h_r_5_34136;
  wire seg_8_4_sp4_h_r_9_34140;
  wire seg_8_4_sp4_r_v_b_12_33895;
  wire seg_8_4_sp4_r_v_b_13_33896;
  wire seg_8_4_sp4_r_v_b_47_34152;
  wire seg_8_4_sp4_v_b_18_30070;
  wire seg_8_5_glb_netwk_0_5;
  wire seg_8_5_glb_netwk_4_9;
  wire seg_8_5_local_g0_2_34160;
  wire seg_8_5_local_g1_1_34167;
  wire seg_8_5_local_g1_5_34171;
  wire seg_8_5_local_g2_5_34179;
  wire seg_8_5_local_g2_7_34181;
  wire seg_8_5_local_g3_3_34185;
  wire seg_8_5_local_g3_4_34186;
  wire seg_8_5_local_g3_5_34187;
  wire seg_8_5_local_g3_7_34189;
  wire seg_8_5_lutff_1_out_30287;
  wire seg_8_5_lutff_3_out_30289;
  wire seg_8_5_lutff_4_out_30290;
  wire seg_8_5_lutff_5_out_30291;
  wire seg_8_5_lutff_7_out_30293;
  wire seg_8_5_sp12_v_b_12_33605;
  wire seg_8_5_sp4_h_l_39_19563;
  wire seg_8_5_sp4_h_r_0_34252;
  wire seg_8_5_sp4_h_r_18_30430;
  wire seg_8_5_sp4_h_r_36_23391;
  wire seg_8_5_sp4_h_r_47_23392;
  wire seg_8_5_sp4_h_r_5_34259;
  wire seg_8_5_sp4_r_v_b_13_34019;
  wire seg_8_5_sp4_v_b_27_30312;
  wire seg_8_5_sp4_v_b_31_30316;
  wire seg_8_5_sp4_v_b_4_30069;
  wire seg_8_5_sp4_v_t_38_30558;
  wire seg_8_5_sp4_v_t_41_30561;
  wire seg_8_5_sp4_v_t_47_30567;
  wire seg_8_6_glb_netwk_0_5;
  wire seg_8_6_glb_netwk_7_12;
  wire seg_8_6_local_g0_3_34284;
  wire seg_8_6_local_g0_5_34286;
  wire seg_8_6_local_g1_5_34294;
  wire seg_8_6_local_g2_1_34298;
  wire seg_8_6_local_g2_3_34300;
  wire seg_8_6_local_g2_7_34304;
  wire seg_8_6_local_g3_1_34306;
  wire seg_8_6_neigh_op_tnr_1_34364;
  wire seg_8_6_sp4_h_l_36_19683;
  wire seg_8_6_sp4_h_l_37_19682;
  wire seg_8_6_sp4_h_l_45_19692;
  wire seg_8_6_sp4_h_r_3_34380;
  wire seg_8_6_sp4_h_r_5_34382;
  wire seg_8_6_sp4_r_v_b_19_34148;
  wire seg_8_6_sp4_r_v_b_29_34268;
  wire seg_8_6_sp4_v_b_22_30320;
  wire seg_8_6_sp4_v_b_26_30436;
  wire seg_8_6_sp4_v_b_30_30440;
  wire seg_8_6_sp4_v_b_31_30439;
  wire seg_8_6_sp4_v_b_32_30442;
  wire seg_8_6_sp4_v_b_33_30441;
  wire seg_8_6_sp4_v_b_35_30443;
  wire seg_8_6_sp4_v_b_3_30189;
  wire seg_8_6_sp4_v_b_40_30560;
  wire seg_8_6_sp4_v_b_44_30564;
  wire seg_8_6_sp4_v_t_37_30680;
  wire seg_8_6_sp4_v_t_47_30690;
  wire seg_8_7_glb_netwk_0_5;
  wire seg_8_7_glb_netwk_5_10;
  wire seg_8_7_local_g0_2_34406;
  wire seg_8_7_local_g0_5_34409;
  wire seg_8_7_local_g1_6_34418;
  wire seg_8_7_sp12_v_b_20_34251;
  wire seg_8_7_sp4_h_l_41_19811;
  wire seg_8_7_sp4_h_l_42_19814;
  wire seg_8_7_sp4_h_l_46_19808;
  wire seg_8_7_sp4_h_r_0_34498;
  wire seg_8_7_sp4_h_r_7_34507;
  wire seg_8_7_sp4_r_v_b_29_34391;
  wire seg_8_7_sp4_v_b_11_30320;
  wire seg_8_7_sp4_v_b_18_30439;
  wire seg_8_7_sp4_v_b_22_30443;
  wire seg_8_7_sp4_v_b_32_30565;
  wire seg_8_7_sp4_v_b_5_30314;
  wire seg_8_7_sp4_v_t_38_30804;
  wire seg_8_7_sp4_v_t_42_30808;
  wire seg_8_8_local_g0_1_34528;
  wire seg_8_8_local_g0_2_34529;
  wire seg_8_8_local_g0_4_34531;
  wire seg_8_8_local_g0_5_34532;
  wire seg_8_8_local_g0_7_34534;
  wire seg_8_8_local_g1_4_34539;
  wire seg_8_8_local_g1_5_34540;
  wire seg_8_8_local_g1_6_34541;
  wire seg_8_8_local_g1_7_34542;
  wire seg_8_8_local_g2_1_34544;
  wire seg_8_8_local_g2_4_34547;
  wire seg_8_8_local_g3_1_34552;
  wire seg_8_8_local_g3_2_34553;
  wire seg_8_8_local_g3_7_34558;
  wire seg_8_8_lutff_1_out_30656;
  wire seg_8_8_lutff_2_out_30657;
  wire seg_8_8_lutff_3_out_30658;
  wire seg_8_8_lutff_4_out_30659;
  wire seg_8_8_lutff_5_out_30660;
  wire seg_8_8_lutff_6_out_30661;
  wire seg_8_8_lutff_7_out_30662;
  wire seg_8_8_neigh_op_bnl_1_27176;
  wire seg_8_8_neigh_op_lft_1_27278;
  wire seg_8_8_neigh_op_lft_2_27279;
  wire seg_8_8_neigh_op_lft_4_27281;
  wire seg_8_8_neigh_op_lft_5_27282;
  wire seg_8_8_neigh_op_lft_6_27283;
  wire seg_8_8_neigh_op_lft_7_27284;
  wire seg_8_8_neigh_op_tnr_1_34610;
  wire seg_8_8_neigh_op_tnr_2_34611;
  wire seg_8_8_neigh_op_tnr_4_34613;
  wire seg_8_8_neigh_op_top_4_30782;
  wire seg_8_8_neigh_op_top_5_30783;
  wire seg_8_8_neigh_op_top_7_30785;
  wire seg_8_8_sp12_v_b_23_34497;
  wire seg_8_8_sp4_h_r_11_34624;
  wire seg_8_8_sp4_h_r_3_34626;
  wire seg_8_8_sp4_h_r_6_34629;
  wire seg_8_8_sp4_h_r_7_34630;
  wire seg_8_8_sp4_h_r_9_34632;
  wire seg_8_8_sp4_v_b_2_30436;
  wire seg_8_8_sp4_v_b_47_30813;
  wire seg_8_8_sp4_v_b_6_30440;
  wire seg_8_8_sp4_v_b_8_30442;
  wire seg_8_8_sp4_v_t_46_30935;
  wire seg_8_9_glb_netwk_0_5;
  wire seg_8_9_glb_netwk_4_9;
  wire seg_8_9_local_g0_2_34652;
  wire seg_8_9_local_g1_4_34662;
  wire seg_8_9_local_g1_6_34664;
  wire seg_8_9_local_g1_7_34665;
  wire seg_8_9_local_g2_2_34668;
  wire seg_8_9_local_g2_6_34672;
  wire seg_8_9_local_g3_2_34676;
  wire seg_8_9_local_g3_4_34678;
  wire seg_8_9_lutff_1_out_30779;
  wire seg_8_9_lutff_2_out_30780;
  wire seg_8_9_lutff_4_out_30782;
  wire seg_8_9_lutff_5_out_30783;
  wire seg_8_9_lutff_6_out_30784;
  wire seg_8_9_lutff_7_out_30785;
  wire seg_8_9_neigh_op_tnl_2_27483;
  wire seg_8_9_neigh_op_tnl_4_27485;
  wire seg_8_9_sp4_h_r_0_34744;
  wire seg_8_9_sp4_h_r_10_34746;
  wire seg_8_9_sp4_h_r_6_34752;
  wire seg_8_9_sp4_r_v_b_1_34387;
  wire seg_8_9_sp4_r_v_b_42_34762;
  wire seg_8_9_sp4_v_b_0_30557;
  wire seg_8_9_sp4_v_b_5_30560;
  wire seg_8_9_sp4_v_b_6_30563;
  wire seg_8_9_sp4_v_b_8_30565;
  wire seg_8_9_sp4_v_b_9_30564;
  wire seg_8_9_sp4_v_t_38_31050;
  wire seg_8_9_sp4_v_t_41_31053;
  wire seg_8_9_sp4_v_t_43_31055;
  wire seg_8_9_sp4_v_t_45_31057;
  wire seg_9_0_local_g0_4_37403;
  wire seg_9_0_local_g0_7_37406;
  wire seg_9_0_span4_horz_r_7_33619;
  wire seg_9_0_span4_vert_20_33749;
  wire seg_9_10_glb_netwk_0_5;
  wire seg_9_10_glb_netwk_4_9;
  wire seg_9_10_local_g0_0_38604;
  wire seg_9_10_local_g0_4_38608;
  wire seg_9_10_local_g1_2_38614;
  wire seg_9_10_local_g1_3_38615;
  wire seg_9_10_local_g1_4_38616;
  wire seg_9_10_local_g2_4_38624;
  wire seg_9_10_local_g3_1_38629;
  wire seg_9_10_local_g3_4_38632;
  wire seg_9_10_lutff_1_out_34733;
  wire seg_9_10_lutff_2_out_34734;
  wire seg_9_10_lutff_4_out_34736;
  wire seg_9_10_lutff_5_out_34737;
  wire seg_9_10_lutff_6_out_34738;
  wire seg_9_10_neigh_op_tnl_4_31028;
  wire seg_9_10_sp4_h_l_38_24010;
  wire seg_9_10_sp4_h_l_41_24011;
  wire seg_9_10_sp4_h_l_42_24014;
  wire seg_9_10_sp4_h_l_43_24013;
  wire seg_9_10_sp4_h_l_44_24016;
  wire seg_9_10_sp4_h_r_11_38701;
  wire seg_9_10_sp4_h_r_19_34875;
  wire seg_9_10_sp4_h_r_2_38702;
  wire seg_9_10_sp4_h_r_3_38703;
  wire seg_9_10_sp4_h_r_8_38708;
  wire seg_9_10_sp4_r_v_b_31_38593;
  wire seg_9_10_sp4_v_b_0_34511;
  wire seg_9_10_sp4_v_b_11_34520;
  wire seg_9_10_sp4_v_b_12_34633;
  wire seg_9_10_sp4_v_b_16_34637;
  wire seg_9_10_sp4_v_b_44_34887;
  wire seg_9_10_sp4_v_b_46_34889;
  wire seg_9_10_sp4_v_t_37_35003;
  wire seg_9_11_glb_netwk_0_5;
  wire seg_9_11_glb_netwk_4_9;
  wire seg_9_11_local_g1_0_38735;
  wire seg_9_11_local_g1_3_38738;
  wire seg_9_11_local_g2_6_38749;
  wire seg_9_11_lutff_0_out_34855;
  wire seg_9_11_lutff_6_out_34861;
  wire seg_9_11_sp4_h_l_39_24132;
  wire seg_9_11_sp4_h_l_40_24135;
  wire seg_9_11_sp4_h_r_12_34991;
  wire seg_9_11_sp4_h_r_16_34997;
  wire seg_9_11_sp4_h_r_28_31165;
  wire seg_9_11_sp4_h_r_32_31169;
  wire seg_9_11_sp4_h_r_44_27738;
  wire seg_9_11_sp4_r_v_b_13_38588;
  wire seg_9_11_sp4_r_v_b_17_38592;
  wire seg_9_11_sp4_r_v_b_1_38464;
  wire seg_9_11_sp4_v_b_0_34634;
  wire seg_9_11_sp4_v_b_12_34756;
  wire seg_9_11_sp4_v_b_16_34760;
  wire seg_9_11_sp4_v_b_19_34763;
  wire seg_9_11_sp4_v_b_28_34884;
  wire seg_9_11_sp4_v_b_2_34636;
  wire seg_9_11_sp4_v_b_44_35010;
  wire seg_9_11_sp4_v_t_38_35127;
  wire seg_9_11_sp4_v_t_42_35131;
  wire seg_9_12_glb_netwk_0_5;
  wire seg_9_12_local_g0_2_38852;
  wire seg_9_12_local_g1_0_38858;
  wire seg_9_12_local_g2_7_38873;
  wire seg_9_12_local_g3_3_38877;
  wire seg_9_12_local_g3_5_38879;
  wire seg_9_12_local_g3_6_38880;
  wire seg_9_12_lutff_5_out_34983;
  wire seg_9_12_neigh_op_bnl_3_31027;
  wire seg_9_12_neigh_op_tnl_5_31275;
  wire seg_9_12_sp12_v_b_1_37438;
  wire seg_9_12_sp4_h_r_0_38944;
  wire seg_9_12_sp4_h_r_16_35120;
  wire seg_9_12_sp4_h_r_18_35122;
  wire seg_9_12_sp4_h_r_2_38948;
  wire seg_9_12_sp4_h_r_9_38955;
  wire seg_9_12_sp4_r_v_b_15_38713;
  wire seg_9_12_sp4_r_v_b_22_38720;
  wire seg_9_12_sp4_v_b_1_34756;
  wire seg_9_12_sp4_v_b_40_35129;
  wire seg_9_12_sp4_v_t_39_35251;
  wire seg_9_12_sp4_v_t_42_35254;
  wire seg_9_13_glb_netwk_0_5;
  wire seg_9_13_local_g1_1_38982;
  wire seg_9_13_local_g1_2_38983;
  wire seg_9_13_local_g1_3_38984;
  wire seg_9_13_local_g2_1_38990;
  wire seg_9_13_local_g2_2_38991;
  wire seg_9_13_local_g3_3_39000;
  wire seg_9_13_local_g3_6_39003;
  wire seg_9_13_lutff_3_out_35104;
  wire seg_9_13_neigh_op_rgt_1_38933;
  wire seg_9_13_sp12_h_r_3_35232;
  wire seg_9_13_sp4_h_r_10_39069;
  wire seg_9_13_sp4_h_r_11_39070;
  wire seg_9_13_sp4_h_r_1_39068;
  wire seg_9_13_sp4_h_r_30_31413;
  wire seg_9_13_sp4_h_r_6_39075;
  wire seg_9_13_sp4_r_v_b_2_38713;
  wire seg_9_13_sp4_r_v_b_34_38967;
  wire seg_9_13_sp4_v_b_11_34889;
  wire seg_9_13_sp4_v_b_28_35130;
  wire seg_9_13_sp4_v_b_4_34884;
  wire seg_9_13_sp4_v_b_5_34883;
  wire seg_9_13_sp4_v_b_7_34885;
  wire seg_9_13_sp4_v_t_37_35372;
  wire seg_9_13_sp4_v_t_39_35374;
  wire seg_9_13_sp4_v_t_43_35378;
  wire seg_9_14_glb_netwk_0_5;
  wire seg_9_14_local_g0_2_39098;
  wire seg_9_14_local_g0_3_39099;
  wire seg_9_14_local_g0_4_39100;
  wire seg_9_14_local_g1_3_39107;
  wire seg_9_14_local_g1_6_39110;
  wire seg_9_14_local_g2_2_39114;
  wire seg_9_14_local_g2_3_39115;
  wire seg_9_14_local_g2_6_39118;
  wire seg_9_14_local_g3_3_39123;
  wire seg_9_14_local_g3_6_39126;
  wire seg_9_14_lutff_0_out_35224;
  wire seg_9_14_lutff_2_out_35226;
  wire seg_9_14_lutff_3_out_35227;
  wire seg_9_14_lutff_4_out_35228;
  wire seg_9_14_lutff_7_out_35231;
  wire seg_9_14_neigh_op_bnr_2_38934;
  wire seg_9_14_sp4_h_r_0_39190;
  wire seg_9_14_sp4_h_r_20_35370;
  wire seg_9_14_sp4_h_r_26_31532;
  wire seg_9_14_sp4_h_r_5_39197;
  wire seg_9_14_sp4_r_v_b_10_38844;
  wire seg_9_14_sp4_r_v_b_19_38963;
  wire seg_9_14_sp4_r_v_b_46_39212;
  wire seg_9_14_sp4_r_v_b_6_38840;
  wire seg_9_14_sp4_v_b_11_35012;
  wire seg_9_14_sp4_v_b_2_35005;
  wire seg_9_14_sp4_v_b_3_35004;
  wire seg_9_14_sp4_v_b_46_35381;
  wire seg_9_14_sp4_v_b_7_35008;
  wire seg_9_14_sp4_v_b_9_35010;
  wire seg_9_14_sp4_v_t_39_35497;
  wire seg_9_14_sp4_v_t_41_35499;
  wire seg_9_15_glb_netwk_0_5;
  wire seg_9_15_local_g0_5_39224;
  wire seg_9_15_local_g1_1_39228;
  wire seg_9_15_local_g1_3_39230;
  wire seg_9_15_local_g1_4_39231;
  wire seg_9_15_local_g1_6_39233;
  wire seg_9_15_local_g1_7_39234;
  wire seg_9_15_local_g2_0_39235;
  wire seg_9_15_local_g2_1_39236;
  wire seg_9_15_local_g2_3_39238;
  wire seg_9_15_local_g3_1_39244;
  wire seg_9_15_local_g3_3_39246;
  wire seg_9_15_local_g3_4_39247;
  wire seg_9_15_local_g3_6_39249;
  wire seg_9_15_lutff_0_out_35347;
  wire seg_9_15_lutff_1_out_35348;
  wire seg_9_15_lutff_3_out_35350;
  wire seg_9_15_lutff_4_out_35351;
  wire seg_9_15_lutff_5_out_35352;
  wire seg_9_15_lutff_6_out_35353;
  wire seg_9_15_lutff_7_out_35354;
  wire seg_9_15_neigh_op_bot_4_35228;
  wire seg_9_15_neigh_op_bot_7_35231;
  wire seg_9_15_neigh_op_rgt_0_39178;
  wire seg_9_15_neigh_op_rgt_4_39182;
  wire seg_9_15_sp12_v_b_9_38327;
  wire seg_9_15_sp4_h_r_21_35492;
  wire seg_9_15_sp4_h_r_27_31656;
  wire seg_9_15_sp4_h_r_36_28136;
  wire seg_9_15_sp4_h_r_3_39318;
  wire seg_9_15_sp4_h_r_4_39319;
  wire seg_9_15_sp4_h_r_6_39321;
  wire seg_9_15_sp4_r_v_b_11_38966;
  wire seg_9_15_sp4_r_v_b_1_38956;
  wire seg_9_15_sp4_r_v_b_22_39089;
  wire seg_9_15_sp4_v_b_25_35371;
  wire seg_9_15_sp4_v_b_2_35128;
  wire seg_9_16_glb_netwk_0_5;
  wire seg_9_16_local_g0_2_39344;
  wire seg_9_16_local_g0_3_39345;
  wire seg_9_16_local_g0_6_39348;
  wire seg_9_16_local_g1_2_39352;
  wire seg_9_16_local_g2_2_39360;
  wire seg_9_16_local_g2_6_39364;
  wire seg_9_16_sp12_h_r_6_28234;
  wire seg_9_16_sp4_h_r_0_39436;
  wire seg_9_16_sp4_h_r_10_39438;
  wire seg_9_16_sp4_h_r_18_35614;
  wire seg_9_16_sp4_r_v_b_14_39204;
  wire seg_9_16_sp4_r_v_b_27_39327;
  wire seg_9_16_sp4_r_v_b_31_39331;
  wire seg_9_16_sp4_r_v_b_41_39453;
  wire seg_9_16_sp4_r_v_b_43_39455;
  wire seg_9_16_sp4_v_b_34_35505;
  wire seg_9_16_sp4_v_b_38_35619;
  wire seg_9_17_glb_netwk_0_5;
  wire seg_9_17_local_g0_1_39466;
  wire seg_9_17_local_g1_1_39474;
  wire seg_9_17_local_g1_3_39476;
  wire seg_9_17_local_g1_7_39480;
  wire seg_9_17_local_g2_0_39481;
  wire seg_9_17_local_g2_1_39482;
  wire seg_9_17_local_g2_2_39483;
  wire seg_9_17_local_g2_3_39484;
  wire seg_9_17_local_g3_3_39492;
  wire seg_9_17_lutff_0_out_35593;
  wire seg_9_17_lutff_2_out_35595;
  wire seg_9_17_lutff_3_out_35596;
  wire seg_9_17_neigh_op_bnr_1_39302;
  wire seg_9_17_neigh_op_bnr_3_39304;
  wire seg_9_17_sp4_h_l_39_24870;
  wire seg_9_17_sp4_r_v_b_11_39212;
  wire seg_9_17_sp4_r_v_b_34_39459;
  wire seg_9_17_sp4_r_v_b_35_39458;
  wire seg_9_17_sp4_r_v_b_9_39210;
  wire seg_9_17_sp4_v_b_1_35371;
  wire seg_9_17_sp4_v_b_23_35505;
  wire seg_9_17_sp4_v_b_7_35377;
  wire seg_9_18_glb_netwk_0_5;
  wire seg_9_18_local_g0_0_39588;
  wire seg_9_18_local_g0_1_39589;
  wire seg_9_18_local_g0_2_39590;
  wire seg_9_18_local_g0_3_39591;
  wire seg_9_18_local_g0_4_39592;
  wire seg_9_18_local_g0_6_39594;
  wire seg_9_18_local_g0_7_39595;
  wire seg_9_18_local_g1_0_39596;
  wire seg_9_18_local_g1_1_39597;
  wire seg_9_18_local_g1_2_39598;
  wire seg_9_18_local_g1_3_39599;
  wire seg_9_18_local_g1_4_39600;
  wire seg_9_18_local_g1_6_39602;
  wire seg_9_18_local_g1_7_39603;
  wire seg_9_18_local_g2_0_39604;
  wire seg_9_18_local_g2_4_39608;
  wire seg_9_18_local_g2_6_39610;
  wire seg_9_18_local_g3_0_39612;
  wire seg_9_18_local_g3_1_39613;
  wire seg_9_18_local_g3_3_39615;
  wire seg_9_18_local_g3_6_39618;
  wire seg_9_18_lutff_0_out_35716;
  wire seg_9_18_lutff_2_out_35718;
  wire seg_9_18_lutff_5_out_35721;
  wire seg_9_18_lutff_6_out_35722;
  wire seg_9_18_lutff_7_out_35723;
  wire seg_9_18_neigh_op_bnr_0_39424;
  wire seg_9_18_neigh_op_bnr_1_39425;
  wire seg_9_18_neigh_op_bnr_2_39426;
  wire seg_9_18_neigh_op_bnr_4_39428;
  wire seg_9_18_neigh_op_bnr_6_39430;
  wire seg_9_18_neigh_op_bnr_7_39431;
  wire seg_9_18_neigh_op_bot_2_35595;
  wire seg_9_18_sp4_h_r_8_39692;
  wire seg_9_18_sp4_r_v_b_12_39448;
  wire seg_9_18_sp4_r_v_b_14_39450;
  wire seg_9_18_sp4_r_v_b_17_39453;
  wire seg_9_18_sp4_r_v_b_19_39455;
  wire seg_9_18_sp4_r_v_b_1_39325;
  wire seg_9_18_sp4_r_v_b_22_39458;
  wire seg_9_18_sp4_r_v_b_27_39573;
  wire seg_9_18_sp4_r_v_b_35_39581;
  wire seg_9_18_sp4_r_v_b_40_39698;
  wire seg_9_18_sp4_r_v_b_4_39330;
  wire seg_9_18_sp4_r_v_b_7_39331;
  wire seg_9_18_sp4_v_b_11_35504;
  wire seg_9_18_sp4_v_b_14_35619;
  wire seg_9_18_sp4_v_b_24_35741;
  wire seg_9_18_sp4_v_b_3_35496;
  wire seg_9_19_sp4_v_b_5_35621;
  wire seg_9_1_glb_netwk_0_5;
  wire seg_9_1_glb_netwk_4_9;
  wire seg_9_1_local_g0_0_37457;
  wire seg_9_1_local_g0_5_37462;
  wire seg_9_1_local_g0_7_37464;
  wire seg_9_1_local_g1_3_37468;
  wire seg_9_1_local_g2_7_37480;
  wire seg_9_1_lutff_1_out_33585;
  wire seg_9_1_lutff_3_out_33587;
  wire seg_9_1_lutff_4_out_33588;
  wire seg_9_1_lutff_6_out_33590;
  wire seg_9_1_lutff_7_out_33591;
  wire seg_9_1_neigh_op_lft_3_29756;
  wire seg_9_1_neigh_op_lft_5_29758;
  wire seg_9_1_neigh_op_lft_7_29760;
  wire seg_9_1_sp4_h_r_4_37561;
  wire seg_9_1_sp4_h_r_8_37565;
  wire seg_9_1_sp4_v_t_37_33896;
  wire seg_9_1_sp4_v_t_39_33898;
  wire seg_9_1_sp4_v_t_45_33904;
  wire seg_9_2_glb_netwk_0_5;
  wire seg_9_2_glb_netwk_3_8;
  wire seg_9_2_local_g1_3_37631;
  wire seg_9_2_local_g1_5_37633;
  wire seg_9_2_lutff_3_out_33715;
  wire seg_9_2_lutff_6_out_33718;
  wire seg_9_2_sp4_h_r_13_33883;
  wire seg_9_2_sp4_h_r_2_37718;
  wire seg_9_2_sp4_h_r_3_37719;
  wire seg_9_2_sp4_v_t_43_34025;
  wire seg_9_3_glb_netwk_0_5;
  wire seg_9_3_local_g0_0_37743;
  wire seg_9_3_local_g0_3_37746;
  wire seg_9_3_local_g0_6_37749;
  wire seg_9_3_local_g1_1_37752;
  wire seg_9_3_local_g1_3_37754;
  wire seg_9_3_local_g2_3_37762;
  wire seg_9_3_lutff_3_out_33874;
  wire seg_9_3_neigh_op_bot_3_33715;
  wire seg_9_3_sp4_h_l_44_23155;
  wire seg_9_3_sp4_h_r_1_37838;
  wire seg_9_3_sp4_h_r_22_34009;
  wire seg_9_3_sp4_h_r_3_37842;
  wire seg_9_3_sp4_h_r_4_37843;
  wire seg_9_3_sp4_h_r_5_37844;
  wire seg_9_3_sp4_h_r_8_37847;
  wire seg_9_3_sp4_v_b_17_33772;
  wire seg_9_3_sp4_v_b_28_33900;
  wire seg_9_3_sp4_v_t_45_34150;
  wire seg_9_3_sp4_v_t_47_34152;
  wire seg_9_4_glb_netwk_0_5;
  wire seg_9_4_local_g0_2_37868;
  wire seg_9_4_local_g0_4_37870;
  wire seg_9_4_local_g0_6_37872;
  wire seg_9_4_local_g0_7_37873;
  wire seg_9_4_local_g1_2_37876;
  wire seg_9_4_local_g1_6_37880;
  wire seg_9_4_local_g2_2_37884;
  wire seg_9_4_local_g2_3_37885;
  wire seg_9_4_local_g3_5_37895;
  wire seg_9_4_lutff_2_out_33996;
  wire seg_9_4_lutff_6_out_34000;
  wire seg_9_4_lutff_7_out_34001;
  wire seg_9_4_neigh_op_rgt_3_37828;
  wire seg_9_4_sp4_h_l_43_23275;
  wire seg_9_4_sp4_h_r_10_37962;
  wire seg_9_4_sp4_h_r_14_34134;
  wire seg_9_4_sp4_h_r_18_34138;
  wire seg_9_4_sp4_h_r_20_34140;
  wire seg_9_4_sp4_h_r_26_30302;
  wire seg_9_4_sp4_h_r_32_30308;
  wire seg_9_4_sp4_h_r_3_37965;
  wire seg_9_4_sp4_h_r_6_37968;
  wire seg_9_4_sp4_r_v_b_31_37855;
  wire seg_9_4_sp4_v_b_45_34150;
  wire seg_9_4_sp4_v_b_5_33771;
  wire seg_9_4_sp4_v_t_36_34264;
  wire seg_9_4_sp4_v_t_40_34268;
  wire seg_9_5_glb_netwk_0_5;
  wire seg_9_5_glb_netwk_4_9;
  wire seg_9_5_local_g0_0_37989;
  wire seg_9_5_local_g0_6_37995;
  wire seg_9_5_local_g1_0_37997;
  wire seg_9_5_local_g1_1_37998;
  wire seg_9_5_local_g2_3_38008;
  wire seg_9_5_local_g2_6_38011;
  wire seg_9_5_local_g3_3_38016;
  wire seg_9_5_lutff_0_out_34117;
  wire seg_9_5_lutff_3_out_34120;
  wire seg_9_5_lutff_6_out_34123;
  wire seg_9_5_sp4_h_l_40_23397;
  wire seg_9_5_sp4_h_r_0_38083;
  wire seg_9_5_sp4_h_r_14_34257;
  wire seg_9_5_sp4_h_r_16_34259;
  wire seg_9_5_sp4_h_r_1_38084;
  wire seg_9_5_sp4_h_r_27_30426;
  wire seg_9_5_sp4_h_r_34_30423;
  wire seg_9_5_sp4_h_r_46_27118;
  wire seg_9_5_sp4_h_r_6_38091;
  wire seg_9_5_sp4_v_b_4_33900;
  wire seg_9_5_sp4_v_b_8_33904;
  wire seg_9_5_sp4_v_t_36_34387;
  wire seg_9_5_sp4_v_t_37_34388;
  wire seg_9_5_sp4_v_t_38_34389;
  wire seg_9_5_sp4_v_t_43_34394;
  wire seg_9_6_glb_netwk_0_5;
  wire seg_9_6_glb_netwk_4_9;
  wire seg_9_6_local_g0_6_38118;
  wire seg_9_6_local_g0_7_38119;
  wire seg_9_6_local_g1_0_38120;
  wire seg_9_6_local_g1_7_38127;
  wire seg_9_6_lutff_0_out_34240;
  wire seg_9_6_lutff_2_out_34242;
  wire seg_9_6_neigh_op_top_7_34370;
  wire seg_9_6_sp4_h_l_37_23513;
  wire seg_9_6_sp4_h_r_0_38206;
  wire seg_9_6_sp4_h_r_22_34378;
  wire seg_9_6_sp4_h_r_5_38213;
  wire seg_9_6_sp4_h_r_6_38214;
  wire seg_9_6_sp4_r_v_b_9_37857;
  wire seg_9_6_sp4_v_b_15_34144;
  wire seg_9_6_sp4_v_t_36_34510;
  wire seg_9_6_sp4_v_t_38_34512;
  wire seg_9_7_glb_netwk_0_5;
  wire seg_9_7_glb_netwk_4_9;
  wire seg_9_7_local_g0_1_38236;
  wire seg_9_7_local_g0_5_38240;
  wire seg_9_7_local_g0_7_38242;
  wire seg_9_7_local_g1_1_38244;
  wire seg_9_7_local_g1_3_38246;
  wire seg_9_7_local_g1_6_38249;
  wire seg_9_7_local_g2_2_38253;
  wire seg_9_7_local_g2_4_38255;
  wire seg_9_7_local_g2_5_38256;
  wire seg_9_7_lutff_0_out_34363;
  wire seg_9_7_lutff_1_out_34364;
  wire seg_9_7_lutff_2_out_34365;
  wire seg_9_7_lutff_3_out_34366;
  wire seg_9_7_lutff_4_out_34367;
  wire seg_9_7_lutff_6_out_34369;
  wire seg_9_7_lutff_7_out_34370;
  wire seg_9_7_neigh_op_top_1_34487;
  wire seg_9_7_sp12_h_r_18_1555;
  wire seg_9_7_sp12_h_r_1_38326;
  wire seg_9_7_sp12_v_b_10_37438;
  wire seg_9_7_sp4_h_r_18_34507;
  wire seg_9_7_sp4_h_r_3_38334;
  wire seg_9_7_sp4_r_v_b_35_38228;
  wire seg_9_7_sp4_r_v_b_3_37974;
  wire seg_9_7_sp4_v_b_17_34269;
  wire seg_9_7_sp4_v_b_23_34275;
  wire seg_9_7_sp4_v_b_37_34511;
  wire seg_9_7_sp4_v_b_5_34145;
  wire seg_9_7_sp4_v_b_6_34148;
  wire seg_9_7_sp4_v_t_37_34634;
  wire seg_9_7_sp4_v_t_43_34640;
  wire seg_9_8_glb_netwk_0_5;
  wire seg_9_8_glb_netwk_4_9;
  wire seg_9_8_local_g0_1_38359;
  wire seg_9_8_local_g0_3_38361;
  wire seg_9_8_local_g0_5_38363;
  wire seg_9_8_local_g0_6_38364;
  wire seg_9_8_local_g0_7_38365;
  wire seg_9_8_local_g1_2_38368;
  wire seg_9_8_local_g1_4_38370;
  wire seg_9_8_local_g1_7_38373;
  wire seg_9_8_local_g2_1_38375;
  wire seg_9_8_local_g2_6_38380;
  wire seg_9_8_lutff_1_out_34487;
  wire seg_9_8_lutff_2_out_34488;
  wire seg_9_8_lutff_3_out_34489;
  wire seg_9_8_lutff_4_out_34490;
  wire seg_9_8_lutff_5_out_34491;
  wire seg_9_8_lutff_6_out_34492;
  wire seg_9_8_neigh_op_lft_1_30656;
  wire seg_9_8_neigh_op_lft_2_30657;
  wire seg_9_8_neigh_op_lft_3_30658;
  wire seg_9_8_neigh_op_lft_4_30659;
  wire seg_9_8_neigh_op_lft_5_30660;
  wire seg_9_8_neigh_op_lft_6_30661;
  wire seg_9_8_neigh_op_lft_7_30662;
  wire seg_9_8_neigh_op_tnl_1_30779;
  wire seg_9_8_sp4_h_l_41_23765;
  wire seg_9_8_sp4_h_l_43_23767;
  wire seg_9_8_sp4_h_l_47_23761;
  wire seg_9_8_sp4_h_r_30_30798;
  wire seg_9_8_sp4_v_b_14_34389;
  wire seg_9_8_sp4_v_b_23_34398;
  wire seg_9_8_sp4_v_b_38_34635;
  wire seg_9_8_sp4_v_t_36_34756;
  wire seg_9_8_sp4_v_t_39_34759;
  wire seg_9_8_sp4_v_t_40_34760;
  wire seg_9_9_glb_netwk_0_5;
  wire seg_9_9_glb_netwk_4_9;
  wire seg_9_9_local_g0_3_38484;
  wire seg_9_9_local_g0_4_38485;
  wire seg_9_9_local_g0_5_38486;
  wire seg_9_9_local_g0_6_38487;
  wire seg_9_9_local_g1_2_38491;
  wire seg_9_9_local_g1_5_38494;
  wire seg_9_9_local_g1_6_38495;
  wire seg_9_9_lutff_0_out_34609;
  wire seg_9_9_lutff_1_out_34610;
  wire seg_9_9_lutff_2_out_34611;
  wire seg_9_9_lutff_3_out_34612;
  wire seg_9_9_lutff_4_out_34613;
  wire seg_9_9_lutff_5_out_34614;
  wire seg_9_9_neigh_op_top_2_34734;
  wire seg_9_9_neigh_op_top_5_34737;
  wire seg_9_9_neigh_op_top_6_34738;
  wire seg_9_9_sp4_h_r_22_34747;
  wire seg_9_9_sp4_v_b_12_34510;
  wire seg_9_9_sp4_v_b_20_34518;
  wire seg_9_9_sp4_v_b_30_34640;
  wire seg_9_9_sp4_v_b_4_34392;
  wire seg_9_9_sp4_v_b_5_34391;
  wire seg_9_9_sp4_v_t_37_34880;
  wire seg_9_9_sp4_v_t_39_34882;
  wire seg_9_9_sp4_v_t_47_34890;
  wire t0;
  wire t1004;
  wire t1013;
  wire t106;
  wire t1083;
  wire t116;
  wire t126;
  wire t146;
  wire t175;
  wire t177;
  wire t178;
  wire t179;
  wire t180;
  wire t181;
  wire t182;
  wire t2;
  wire t207;
  wire t209;
  wire t210;
  wire t211;
  wire t212;
  wire t213;
  wire t214;
  wire t264;
  wire t270;
  wire t3;
  wire t36;
  wire t371;
  wire t379;
  wire t383;
  wire t404;
  wire t41;
  wire t412;
  wire t414;
  wire t415;
  wire t416;
  wire t417;
  wire t418;
  wire t419;
  wire t442;
  wire t445;
  wire t447;
  wire t449;
  wire t451;
  wire t453;
  wire t455;
  wire t46;
  wire t471;
  wire t5;
  wire t501;
  wire t549;
  wire t552;
  wire t558;
  wire t591;
  wire t593;
  wire t636;
  wire t638;
  wire t650;
  wire t653;
  wire t654;
  wire t655;
  wire t686;
  wire t688;
  wire t744;
  wire t746;
  wire t784;
  wire t786;
  wire t791;
  wire t802;
  wire t804;
  wire t826;
  wire t835;
  wire t85;
  wire t853;
  wire t862;
  wire t867;
  wire t917;
  wire t929;
  wire t94;
  wire t948;
  wire t957;
  wire t968;
  wire t980;
  wire t987;
  assign net_10 = seg_17_2_glb_netwk_5_10;
  assign net_10015 = seg_1_23_local_g3_2_10015;
  assign net_100150 = seg_25_11_local_g0_0_100150;
  assign net_100154 = seg_25_11_local_g0_4_100154;
  assign net_100155 = seg_25_11_local_g0_5_100155;
  assign net_100156 = seg_25_11_local_g0_6_100156;
  assign net_100164 = seg_25_11_local_g1_6_100164;
  assign net_100168 = seg_25_11_local_g2_2_100168;
  assign net_100169 = seg_25_11_local_g2_3_100169;
  assign net_100170 = seg_25_11_local_g2_4_100170;
  assign net_100171 = seg_25_11_local_g2_5_100171;
  assign net_100172 = seg_25_11_local_g2_6_100172;
  assign net_100173 = seg_25_11_local_g2_7_100173;
  assign net_100175 = seg_25_11_local_g3_1_100175;
  assign net_100176 = seg_25_11_local_g3_2_100176;
  assign net_100178 = seg_25_11_local_g3_4_100178;
  assign net_100180 = seg_25_11_local_g3_6_100180;
  assign net_100181 = seg_25_11_local_g3_7_100181;
  assign net_100302 = seg_25_12_local_g0_2_100302;
  assign net_100303 = seg_25_12_local_g0_3_100303;
  assign net_100309 = seg_25_12_local_g1_1_100309;
  assign net_100310 = seg_25_12_local_g1_2_100310;
  assign net_100311 = seg_25_12_local_g1_3_100311;
  assign net_100312 = seg_25_12_local_g1_4_100312;
  assign net_100313 = seg_25_12_local_g1_5_100313;
  assign net_100314 = seg_25_12_local_g1_6_100314;
  assign net_100317 = seg_25_12_local_g2_1_100317;
  assign net_100318 = seg_25_12_local_g2_2_100318;
  assign net_100319 = seg_25_12_local_g2_3_100319;
  assign net_100320 = seg_25_12_local_g2_4_100320;
  assign net_100325 = seg_25_12_local_g3_1_100325;
  assign net_100326 = seg_25_12_local_g3_2_100326;
  assign net_100330 = seg_25_12_local_g3_6_100330;
  assign net_100331 = seg_25_12_local_g3_7_100331;
  assign net_11272 = seg_2_1_local_g0_1_11272;
  assign net_11278 = seg_2_1_local_g0_7_11278;
  assign net_11279 = seg_2_1_local_g1_0_11279;
  assign net_11283 = seg_2_1_local_g1_4_11283;
  assign net_11293 = seg_2_1_local_g2_6_11293;
  assign net_11294 = seg_2_1_local_g2_7_11294;
  assign net_11295 = seg_2_1_local_g3_0_11295;
  assign net_11302 = seg_2_1_local_g3_7_11302;
  assign net_11435 = seg_2_2_local_g0_1_11435;
  assign net_11436 = seg_2_2_local_g0_2_11436;
  assign net_11437 = seg_2_2_local_g0_3_11437;
  assign net_11438 = seg_2_2_local_g0_4_11438;
  assign net_11439 = seg_2_2_local_g0_5_11439;
  assign net_11440 = seg_2_2_local_g0_6_11440;
  assign net_11442 = seg_2_2_local_g1_0_11442;
  assign net_11444 = seg_2_2_local_g1_2_11444;
  assign net_11445 = seg_2_2_local_g1_3_11445;
  assign net_11446 = seg_2_2_local_g1_4_11446;
  assign net_11447 = seg_2_2_local_g1_5_11447;
  assign net_11448 = seg_2_2_local_g1_6_11448;
  assign net_11449 = seg_2_2_local_g1_7_11449;
  assign net_11451 = seg_2_2_local_g2_1_11451;
  assign net_11452 = seg_2_2_local_g2_2_11452;
  assign net_11454 = seg_2_2_local_g2_4_11454;
  assign net_11455 = seg_2_2_local_g2_5_11455;
  assign net_11462 = seg_2_2_local_g3_4_11462;
  assign net_11465 = seg_2_2_local_g3_7_11465;
  assign net_11558 = seg_2_3_local_g0_1_11558;
  assign net_11560 = seg_2_3_local_g0_3_11560;
  assign net_11561 = seg_2_3_local_g0_4_11561;
  assign net_11562 = seg_2_3_local_g0_5_11562;
  assign net_11563 = seg_2_3_local_g0_6_11563;
  assign net_11564 = seg_2_3_local_g0_7_11564;
  assign net_11565 = seg_2_3_local_g1_0_11565;
  assign net_11567 = seg_2_3_local_g1_2_11567;
  assign net_11569 = seg_2_3_local_g1_4_11569;
  assign net_11570 = seg_2_3_local_g1_5_11570;
  assign net_11572 = seg_2_3_local_g1_7_11572;
  assign net_11573 = seg_2_3_local_g2_0_11573;
  assign net_11575 = seg_2_3_local_g2_2_11575;
  assign net_11585 = seg_2_3_local_g3_4_11585;
  assign net_11586 = seg_2_3_local_g3_5_11586;
  assign net_11588 = seg_2_3_local_g3_7_11588;
  assign net_11680 = seg_2_4_local_g0_0_11680;
  assign net_11682 = seg_2_4_local_g0_2_11682;
  assign net_11683 = seg_2_4_local_g0_3_11683;
  assign net_11684 = seg_2_4_local_g0_4_11684;
  assign net_11686 = seg_2_4_local_g0_6_11686;
  assign net_11690 = seg_2_4_local_g1_2_11690;
  assign net_11692 = seg_2_4_local_g1_4_11692;
  assign net_11693 = seg_2_4_local_g1_5_11693;
  assign net_11695 = seg_2_4_local_g1_7_11695;
  assign net_11696 = seg_2_4_local_g2_0_11696;
  assign net_11699 = seg_2_4_local_g2_3_11699;
  assign net_11702 = seg_2_4_local_g2_6_11702;
  assign net_11704 = seg_2_4_local_g3_0_11704;
  assign net_11706 = seg_2_4_local_g3_2_11706;
  assign net_11707 = seg_2_4_local_g3_3_11707;
  assign net_11708 = seg_2_4_local_g3_4_11708;
  assign net_11709 = seg_2_4_local_g3_5_11709;
  assign net_11710 = seg_2_4_local_g3_6_11710;
  assign net_11809 = seg_2_5_local_g0_6_11809;
  assign net_11816 = seg_2_5_local_g1_5_11816;
  assign net_11819 = seg_2_5_local_g2_0_11819;
  assign net_11821 = seg_2_5_local_g2_2_11821;
  assign net_11825 = seg_2_5_local_g2_6_11825;
  assign net_11829 = seg_2_5_local_g3_2_11829;
  assign net_11831 = seg_2_5_local_g3_4_11831;
  assign net_11833 = seg_2_5_local_g3_6_11833;
  assign net_11930 = seg_2_6_local_g0_4_11930;
  assign net_11941 = seg_2_6_local_g1_7_11941;
  assign net_11943 = seg_2_6_local_g2_1_11943;
  assign net_11950 = seg_2_6_local_g3_0_11950;
  assign net_11954 = seg_2_6_local_g3_4_11954;
  assign net_11956 = seg_2_6_local_g3_6_11956;
  assign net_11957 = seg_2_6_local_g3_7_11957;
  assign net_12 = seg_15_2_glb_netwk_7_12;
  assign net_12050 = seg_2_7_local_g0_1_12050;
  assign net_12053 = seg_2_7_local_g0_4_12053;
  assign net_12054 = seg_2_7_local_g0_5_12054;
  assign net_12056 = seg_2_7_local_g0_7_12056;
  assign net_12065 = seg_2_7_local_g2_0_12065;
  assign net_12067 = seg_2_7_local_g2_2_12067;
  assign net_12071 = seg_2_7_local_g2_6_12071;
  assign net_12073 = seg_2_7_local_g3_0_12073;
  assign net_12077 = seg_2_7_local_g3_4_12077;
  assign net_12172 = seg_2_8_local_g0_0_12172;
  assign net_12174 = seg_2_8_local_g0_2_12174;
  assign net_12175 = seg_2_8_local_g0_3_12175;
  assign net_12176 = seg_2_8_local_g0_4_12176;
  assign net_12177 = seg_2_8_local_g0_5_12177;
  assign net_12178 = seg_2_8_local_g0_6_12178;
  assign net_12179 = seg_2_8_local_g0_7_12179;
  assign net_12180 = seg_2_8_local_g1_0_12180;
  assign net_12181 = seg_2_8_local_g1_1_12181;
  assign net_12182 = seg_2_8_local_g1_2_12182;
  assign net_12183 = seg_2_8_local_g1_3_12183;
  assign net_12184 = seg_2_8_local_g1_4_12184;
  assign net_12186 = seg_2_8_local_g1_6_12186;
  assign net_12187 = seg_2_8_local_g1_7_12187;
  assign net_12190 = seg_2_8_local_g2_2_12190;
  assign net_12193 = seg_2_8_local_g2_5_12193;
  assign net_12194 = seg_2_8_local_g2_6_12194;
  assign net_12201 = seg_2_8_local_g3_5_12201;
  assign net_12295 = seg_2_9_local_g0_0_12295;
  assign net_12297 = seg_2_9_local_g0_2_12297;
  assign net_12299 = seg_2_9_local_g0_4_12299;
  assign net_12300 = seg_2_9_local_g0_5_12300;
  assign net_12302 = seg_2_9_local_g0_7_12302;
  assign net_12308 = seg_2_9_local_g1_5_12308;
  assign net_12312 = seg_2_9_local_g2_1_12312;
  assign net_12319 = seg_2_9_local_g3_0_12319;
  assign net_12419 = seg_2_10_local_g0_1_12419;
  assign net_12432 = seg_2_10_local_g1_6_12432;
  assign net_12433 = seg_2_10_local_g1_7_12433;
  assign net_12436 = seg_2_10_local_g2_2_12436;
  assign net_12439 = seg_2_10_local_g2_5_12439;
  assign net_12442 = seg_2_10_local_g3_0_12442;
  assign net_12443 = seg_2_10_local_g3_1_12443;
  assign net_12446 = seg_2_10_local_g3_4_12446;
  assign net_12541 = seg_2_11_local_g0_0_12541;
  assign net_12542 = seg_2_11_local_g0_1_12542;
  assign net_12544 = seg_2_11_local_g0_3_12544;
  assign net_12546 = seg_2_11_local_g0_5_12546;
  assign net_12553 = seg_2_11_local_g1_4_12553;
  assign net_12554 = seg_2_11_local_g1_5_12554;
  assign net_12556 = seg_2_11_local_g1_7_12556;
  assign net_12559 = seg_2_11_local_g2_2_12559;
  assign net_12563 = seg_2_11_local_g2_6_12563;
  assign net_12564 = seg_2_11_local_g2_7_12564;
  assign net_12565 = seg_2_11_local_g3_0_12565;
  assign net_12566 = seg_2_11_local_g3_1_12566;
  assign net_12567 = seg_2_11_local_g3_2_12567;
  assign net_12568 = seg_2_11_local_g3_3_12568;
  assign net_12569 = seg_2_11_local_g3_4_12569;
  assign net_1257 = seg_0_6_local_g0_3_1257;
  assign net_12570 = seg_2_11_local_g3_5_12570;
  assign net_1258 = seg_0_6_local_g0_4_1258;
  assign net_1259 = seg_0_6_local_g0_5_1259;
  assign net_1262 = seg_0_6_local_g1_0_1262;
  assign net_1264 = seg_0_6_local_g1_2_1264;
  assign net_12667 = seg_2_12_local_g0_3_12667;
  assign net_12669 = seg_2_12_local_g0_5_12669;
  assign net_1267 = seg_0_6_local_g1_5_1267;
  assign net_1268 = seg_0_6_local_g1_6_1268;
  assign net_12681 = seg_2_12_local_g2_1_12681;
  assign net_12683 = seg_2_12_local_g2_3_12683;
  assign net_12685 = seg_2_12_local_g2_5_12685;
  assign net_12688 = seg_2_12_local_g3_0_12688;
  assign net_12690 = seg_2_12_local_g3_2_12690;
  assign net_12692 = seg_2_12_local_g3_4_12692;
  assign net_12695 = seg_2_12_local_g3_7_12695;
  assign net_1272 = seg_0_6_local_g2_2_1272;
  assign net_1274 = seg_0_6_local_g2_4_1274;
  assign net_1275 = seg_0_6_local_g2_5_1275;
  assign net_1276 = seg_0_6_local_g2_6_1276;
  assign net_1278 = seg_0_6_local_g3_0_1278;
  assign net_1279 = seg_0_6_local_g3_1_1279;
  assign net_12790 = seg_2_13_local_g0_3_12790;
  assign net_12793 = seg_2_13_local_g0_6_12793;
  assign net_12798 = seg_2_13_local_g1_3_12798;
  assign net_1280 = seg_0_6_local_g3_2_1280;
  assign net_12802 = seg_2_13_local_g1_7_12802;
  assign net_12804 = seg_2_13_local_g2_1_12804;
  assign net_1281 = seg_0_6_local_g3_3_1281;
  assign net_12810 = seg_2_13_local_g2_7_12810;
  assign net_12812 = seg_2_13_local_g3_1_12812;
  assign net_12814 = seg_2_13_local_g3_3_12814;
  assign net_12816 = seg_2_13_local_g3_5_12816;
  assign net_12818 = seg_2_13_local_g3_7_12818;
  assign net_1285 = seg_0_6_local_g3_7_1285;
  assign net_12913 = seg_2_14_local_g0_3_12913;
  assign net_12919 = seg_2_14_local_g1_1_12919;
  assign net_12920 = seg_2_14_local_g1_2_12920;
  assign net_12925 = seg_2_14_local_g1_7_12925;
  assign net_12927 = seg_2_14_local_g2_1_12927;
  assign net_12928 = seg_2_14_local_g2_2_12928;
  assign net_12931 = seg_2_14_local_g2_5_12931;
  assign net_12932 = seg_2_14_local_g2_6_12932;
  assign net_12934 = seg_2_14_local_g3_0_12934;
  assign net_12935 = seg_2_14_local_g3_1_12935;
  assign net_13034 = seg_2_15_local_g0_1_13034;
  assign net_13035 = seg_2_15_local_g0_2_13035;
  assign net_13036 = seg_2_15_local_g0_3_13036;
  assign net_13037 = seg_2_15_local_g0_4_13037;
  assign net_13039 = seg_2_15_local_g0_6_13039;
  assign net_13040 = seg_2_15_local_g0_7_13040;
  assign net_13043 = seg_2_15_local_g1_2_13043;
  assign net_13055 = seg_2_15_local_g2_6_13055;
  assign net_13060 = seg_2_15_local_g3_3_13060;
  assign net_13062 = seg_2_15_local_g3_5_13062;
  assign net_13063 = seg_2_15_local_g3_6_13063;
  assign net_13158 = seg_2_16_local_g0_2_13158;
  assign net_13163 = seg_2_16_local_g0_7_13163;
  assign net_13164 = seg_2_16_local_g1_0_13164;
  assign net_13166 = seg_2_16_local_g1_2_13166;
  assign net_13173 = seg_2_16_local_g2_1_13173;
  assign net_13174 = seg_2_16_local_g2_2_13174;
  assign net_13183 = seg_2_16_local_g3_3_13183;
  assign net_13187 = seg_2_16_local_g3_7_13187;
  assign net_13291 = seg_2_17_local_g1_4_13291;
  assign net_13294 = seg_2_17_local_g1_7_13294;
  assign net_13301 = seg_2_17_local_g2_6_13301;
  assign net_13403 = seg_2_18_local_g0_1_13403;
  assign net_13407 = seg_2_18_local_g0_5_13407;
  assign net_13408 = seg_2_18_local_g0_6_13408;
  assign net_13409 = seg_2_18_local_g0_7_13409;
  assign net_13421 = seg_2_18_local_g2_3_13421;
  assign net_13528 = seg_2_19_local_g0_3_13528;
  assign net_13529 = seg_2_19_local_g0_4_13529;
  assign net_13531 = seg_2_19_local_g0_6_13531;
  assign net_13533 = seg_2_19_local_g1_0_13533;
  assign net_13537 = seg_2_19_local_g1_4_13537;
  assign net_13538 = seg_2_19_local_g1_5_13538;
  assign net_13540 = seg_2_19_local_g1_7_13540;
  assign net_13650 = seg_2_20_local_g0_2_13650;
  assign net_13652 = seg_2_20_local_g0_4_13652;
  assign net_13653 = seg_2_20_local_g0_5_13653;
  assign net_13655 = seg_2_20_local_g0_7_13655;
  assign net_13672 = seg_2_20_local_g3_0_13672;
  assign net_13776 = seg_2_21_local_g0_5_13776;
  assign net_13779 = seg_2_21_local_g1_0_13779;
  assign net_13897 = seg_2_22_local_g0_3_13897;
  assign net_13920 = seg_2_22_local_g3_2_13920;
  assign net_14026 = seg_2_23_local_g1_1_14026;
  assign net_1461 = seg_0_7_local_g0_1_1461;
  assign net_1464 = seg_0_7_local_g0_4_1464;
  assign net_1471 = seg_0_7_local_g1_3_1471;
  assign net_1474 = seg_0_7_local_g1_6_1474;
  assign net_1476 = seg_0_7_local_g2_0_1476;
  assign net_1478 = seg_0_7_local_g2_2_1478;
  assign net_1479 = seg_0_7_local_g2_3_1479;
  assign net_1483 = seg_0_7_local_g2_7_1483;
  assign net_1484 = seg_0_7_local_g3_0_1484;
  assign net_1485 = seg_0_7_local_g3_1_1485;
  assign net_1486 = seg_0_7_local_g3_2_1486;
  assign net_1487 = seg_0_7_local_g3_3_1487;
  assign net_1488 = seg_0_7_local_g3_4_1488;
  assign net_1489 = seg_0_7_local_g3_5_1489;
  assign net_1490 = seg_0_7_local_g3_6_1490;
  assign net_1491 = seg_0_7_local_g3_7_1491;
  assign net_15103 = seg_3_1_local_g0_1_15103;
  assign net_15104 = seg_3_1_local_g0_2_15104;
  assign net_15106 = seg_3_1_local_g0_4_15106;
  assign net_15110 = seg_3_1_local_g1_0_15110;
  assign net_15115 = seg_3_1_local_g1_5_15115;
  assign net_15118 = seg_3_1_local_g2_0_15118;
  assign net_15119 = seg_3_1_local_g2_1_15119;
  assign net_15120 = seg_3_1_local_g2_2_15120;
  assign net_15121 = seg_3_1_local_g2_3_15121;
  assign net_15122 = seg_3_1_local_g2_4_15122;
  assign net_15124 = seg_3_1_local_g2_6_15124;
  assign net_15126 = seg_3_1_local_g3_0_15126;
  assign net_15127 = seg_3_1_local_g3_1_15127;
  assign net_15129 = seg_3_1_local_g3_3_15129;
  assign net_15131 = seg_3_1_local_g3_5_15131;
  assign net_15132 = seg_3_1_local_g3_6_15132;
  assign net_15133 = seg_3_1_local_g3_7_15133;
  assign net_15265 = seg_3_2_local_g0_0_15265;
  assign net_15268 = seg_3_2_local_g0_3_15268;
  assign net_15269 = seg_3_2_local_g0_4_15269;
  assign net_15270 = seg_3_2_local_g0_5_15270;
  assign net_15273 = seg_3_2_local_g1_0_15273;
  assign net_15274 = seg_3_2_local_g1_1_15274;
  assign net_15279 = seg_3_2_local_g1_6_15279;
  assign net_15280 = seg_3_2_local_g1_7_15280;
  assign net_15282 = seg_3_2_local_g2_1_15282;
  assign net_15283 = seg_3_2_local_g2_2_15283;
  assign net_15284 = seg_3_2_local_g2_3_15284;
  assign net_15285 = seg_3_2_local_g2_4_15285;
  assign net_15286 = seg_3_2_local_g2_5_15286;
  assign net_15289 = seg_3_2_local_g3_0_15289;
  assign net_15290 = seg_3_2_local_g3_1_15290;
  assign net_15291 = seg_3_2_local_g3_2_15291;
  assign net_15292 = seg_3_2_local_g3_3_15292;
  assign net_15293 = seg_3_2_local_g3_4_15293;
  assign net_15294 = seg_3_2_local_g3_5_15294;
  assign net_15295 = seg_3_2_local_g3_6_15295;
  assign net_15296 = seg_3_2_local_g3_7_15296;
  assign net_15390 = seg_3_3_local_g0_2_15390;
  assign net_15391 = seg_3_3_local_g0_3_15391;
  assign net_15392 = seg_3_3_local_g0_4_15392;
  assign net_15394 = seg_3_3_local_g0_6_15394;
  assign net_15395 = seg_3_3_local_g0_7_15395;
  assign net_15397 = seg_3_3_local_g1_1_15397;
  assign net_15398 = seg_3_3_local_g1_2_15398;
  assign net_15399 = seg_3_3_local_g1_3_15399;
  assign net_15400 = seg_3_3_local_g1_4_15400;
  assign net_15402 = seg_3_3_local_g1_6_15402;
  assign net_15404 = seg_3_3_local_g2_0_15404;
  assign net_15406 = seg_3_3_local_g2_2_15406;
  assign net_15407 = seg_3_3_local_g2_3_15407;
  assign net_15408 = seg_3_3_local_g2_4_15408;
  assign net_15409 = seg_3_3_local_g2_5_15409;
  assign net_15410 = seg_3_3_local_g2_6_15410;
  assign net_15412 = seg_3_3_local_g3_0_15412;
  assign net_15414 = seg_3_3_local_g3_2_15414;
  assign net_15415 = seg_3_3_local_g3_3_15415;
  assign net_15416 = seg_3_3_local_g3_4_15416;
  assign net_15417 = seg_3_3_local_g3_5_15417;
  assign net_15511 = seg_3_4_local_g0_0_15511;
  assign net_15514 = seg_3_4_local_g0_3_15514;
  assign net_15516 = seg_3_4_local_g0_5_15516;
  assign net_15518 = seg_3_4_local_g0_7_15518;
  assign net_15519 = seg_3_4_local_g1_0_15519;
  assign net_15522 = seg_3_4_local_g1_3_15522;
  assign net_15523 = seg_3_4_local_g1_4_15523;
  assign net_15524 = seg_3_4_local_g1_5_15524;
  assign net_15525 = seg_3_4_local_g1_6_15525;
  assign net_15526 = seg_3_4_local_g1_7_15526;
  assign net_15527 = seg_3_4_local_g2_0_15527;
  assign net_15530 = seg_3_4_local_g2_3_15530;
  assign net_15533 = seg_3_4_local_g2_6_15533;
  assign net_15536 = seg_3_4_local_g3_1_15536;
  assign net_15638 = seg_3_5_local_g0_4_15638;
  assign net_15640 = seg_3_5_local_g0_6_15640;
  assign net_15642 = seg_3_5_local_g1_0_15642;
  assign net_15644 = seg_3_5_local_g1_2_15644;
  assign net_15648 = seg_3_5_local_g1_6_15648;
  assign net_15651 = seg_3_5_local_g2_1_15651;
  assign net_15653 = seg_3_5_local_g2_3_15653;
  assign net_15655 = seg_3_5_local_g2_5_15655;
  assign net_15660 = seg_3_5_local_g3_2_15660;
  assign net_15761 = seg_3_6_local_g0_4_15761;
  assign net_15762 = seg_3_6_local_g0_5_15762;
  assign net_15765 = seg_3_6_local_g1_0_15765;
  assign net_15766 = seg_3_6_local_g1_1_15766;
  assign net_15767 = seg_3_6_local_g1_2_15767;
  assign net_15770 = seg_3_6_local_g1_5_15770;
  assign net_15772 = seg_3_6_local_g1_7_15772;
  assign net_15774 = seg_3_6_local_g2_1_15774;
  assign net_15775 = seg_3_6_local_g2_2_15775;
  assign net_15776 = seg_3_6_local_g2_3_15776;
  assign net_15781 = seg_3_6_local_g3_0_15781;
  assign net_15783 = seg_3_6_local_g3_2_15783;
  assign net_15784 = seg_3_6_local_g3_3_15784;
  assign net_15882 = seg_3_7_local_g0_2_15882;
  assign net_15883 = seg_3_7_local_g0_3_15883;
  assign net_15884 = seg_3_7_local_g0_4_15884;
  assign net_15885 = seg_3_7_local_g0_5_15885;
  assign net_15886 = seg_3_7_local_g0_6_15886;
  assign net_15888 = seg_3_7_local_g1_0_15888;
  assign net_15889 = seg_3_7_local_g1_1_15889;
  assign net_15890 = seg_3_7_local_g1_2_15890;
  assign net_15891 = seg_3_7_local_g1_3_15891;
  assign net_15892 = seg_3_7_local_g1_4_15892;
  assign net_15894 = seg_3_7_local_g1_6_15894;
  assign net_15895 = seg_3_7_local_g1_7_15895;
  assign net_16003 = seg_3_8_local_g0_0_16003;
  assign net_16005 = seg_3_8_local_g0_2_16005;
  assign net_16013 = seg_3_8_local_g1_2_16013;
  assign net_16020 = seg_3_8_local_g2_1_16020;
  assign net_16023 = seg_3_8_local_g2_4_16023;
  assign net_16029 = seg_3_8_local_g3_2_16029;
  assign net_16127 = seg_3_9_local_g0_1_16127;
  assign net_16129 = seg_3_9_local_g0_3_16129;
  assign net_16130 = seg_3_9_local_g0_4_16130;
  assign net_16132 = seg_3_9_local_g0_6_16132;
  assign net_16133 = seg_3_9_local_g0_7_16133;
  assign net_16134 = seg_3_9_local_g1_0_16134;
  assign net_16135 = seg_3_9_local_g1_1_16135;
  assign net_16138 = seg_3_9_local_g1_4_16138;
  assign net_16139 = seg_3_9_local_g1_5_16139;
  assign net_16141 = seg_3_9_local_g1_7_16141;
  assign net_16142 = seg_3_9_local_g2_0_16142;
  assign net_16149 = seg_3_9_local_g2_7_16149;
  assign net_16153 = seg_3_9_local_g3_3_16153;
  assign net_16156 = seg_3_9_local_g3_6_16156;
  assign net_16253 = seg_3_10_local_g0_4_16253;
  assign net_16254 = seg_3_10_local_g0_5_16254;
  assign net_16260 = seg_3_10_local_g1_3_16260;
  assign net_16261 = seg_3_10_local_g1_4_16261;
  assign net_16268 = seg_3_10_local_g2_3_16268;
  assign net_16273 = seg_3_10_local_g3_0_16273;
  assign net_16276 = seg_3_10_local_g3_3_16276;
  assign net_16278 = seg_3_10_local_g3_5_16278;
  assign net_16375 = seg_3_11_local_g0_3_16375;
  assign net_16383 = seg_3_11_local_g1_3_16383;
  assign net_16385 = seg_3_11_local_g1_5_16385;
  assign net_16386 = seg_3_11_local_g1_6_16386;
  assign net_16387 = seg_3_11_local_g1_7_16387;
  assign net_16388 = seg_3_11_local_g2_0_16388;
  assign net_16390 = seg_3_11_local_g2_2_16390;
  assign net_16394 = seg_3_11_local_g2_6_16394;
  assign net_16498 = seg_3_12_local_g0_3_16498;
  assign net_16499 = seg_3_12_local_g0_4_16499;
  assign net_16500 = seg_3_12_local_g0_5_16500;
  assign net_16504 = seg_3_12_local_g1_1_16504;
  assign net_16507 = seg_3_12_local_g1_4_16507;
  assign net_16508 = seg_3_12_local_g1_5_16508;
  assign net_16510 = seg_3_12_local_g1_7_16510;
  assign net_16513 = seg_3_12_local_g2_2_16513;
  assign net_16514 = seg_3_12_local_g2_3_16514;
  assign net_16515 = seg_3_12_local_g2_4_16515;
  assign net_16517 = seg_3_12_local_g2_6_16517;
  assign net_16518 = seg_3_12_local_g2_7_16518;
  assign net_16523 = seg_3_12_local_g3_4_16523;
  assign net_16525 = seg_3_12_local_g3_6_16525;
  assign net_16623 = seg_3_13_local_g0_5_16623;
  assign net_16625 = seg_3_13_local_g0_7_16625;
  assign net_16633 = seg_3_13_local_g1_7_16633;
  assign net_16634 = seg_3_13_local_g2_0_16634;
  assign net_16636 = seg_3_13_local_g2_2_16636;
  assign net_16637 = seg_3_13_local_g2_3_16637;
  assign net_16638 = seg_3_13_local_g2_4_16638;
  assign net_16639 = seg_3_13_local_g2_5_16639;
  assign net_16640 = seg_3_13_local_g2_6_16640;
  assign net_16642 = seg_3_13_local_g3_0_16642;
  assign net_16643 = seg_3_13_local_g3_1_16643;
  assign net_16644 = seg_3_13_local_g3_2_16644;
  assign net_16645 = seg_3_13_local_g3_3_16645;
  assign net_16646 = seg_3_13_local_g3_4_16646;
  assign net_16647 = seg_3_13_local_g3_5_16647;
  assign net_16648 = seg_3_13_local_g3_6_16648;
  assign net_16742 = seg_3_14_local_g0_1_16742;
  assign net_16748 = seg_3_14_local_g0_7_16748;
  assign net_16756 = seg_3_14_local_g1_7_16756;
  assign net_16757 = seg_3_14_local_g2_0_16757;
  assign net_16758 = seg_3_14_local_g2_1_16758;
  assign net_16761 = seg_3_14_local_g2_4_16761;
  assign net_16762 = seg_3_14_local_g2_5_16762;
  assign net_16765 = seg_3_14_local_g3_0_16765;
  assign net_16767 = seg_3_14_local_g3_2_16767;
  assign net_16768 = seg_3_14_local_g3_3_16768;
  assign net_16770 = seg_3_14_local_g3_5_16770;
  assign net_16864 = seg_3_15_local_g0_0_16864;
  assign net_16866 = seg_3_15_local_g0_2_16866;
  assign net_16867 = seg_3_15_local_g0_3_16867;
  assign net_16868 = seg_3_15_local_g0_4_16868;
  assign net_16869 = seg_3_15_local_g0_5_16869;
  assign net_16873 = seg_3_15_local_g1_1_16873;
  assign net_16878 = seg_3_15_local_g1_6_16878;
  assign net_16883 = seg_3_15_local_g2_3_16883;
  assign net_16884 = seg_3_15_local_g2_4_16884;
  assign net_16886 = seg_3_15_local_g2_6_16886;
  assign net_16890 = seg_3_15_local_g3_2_16890;
  assign net_16892 = seg_3_15_local_g3_4_16892;
  assign net_16893 = seg_3_15_local_g3_5_16893;
  assign net_16894 = seg_3_15_local_g3_6_16894;
  assign net_16989 = seg_3_16_local_g0_2_16989;
  assign net_16990 = seg_3_16_local_g0_3_16990;
  assign net_16992 = seg_3_16_local_g0_5_16992;
  assign net_16998 = seg_3_16_local_g1_3_16998;
  assign net_16999 = seg_3_16_local_g1_4_16999;
  assign net_17001 = seg_3_16_local_g1_6_17001;
  assign net_17004 = seg_3_16_local_g2_1_17004;
  assign net_17016 = seg_3_16_local_g3_5_17016;
  assign net_17114 = seg_3_17_local_g0_4_17114;
  assign net_17115 = seg_3_17_local_g0_5_17115;
  assign net_17121 = seg_3_17_local_g1_3_17121;
  assign net_17126 = seg_3_17_local_g2_0_17126;
  assign net_17127 = seg_3_17_local_g2_1_17127;
  assign net_17132 = seg_3_17_local_g2_6_17132;
  assign net_17133 = seg_3_17_local_g2_7_17133;
  assign net_17233 = seg_3_18_local_g0_0_17233;
  assign net_17234 = seg_3_18_local_g0_1_17234;
  assign net_17237 = seg_3_18_local_g0_4_17237;
  assign net_17238 = seg_3_18_local_g0_5_17238;
  assign net_17241 = seg_3_18_local_g1_0_17241;
  assign net_17242 = seg_3_18_local_g1_1_17242;
  assign net_17243 = seg_3_18_local_g1_2_17243;
  assign net_17244 = seg_3_18_local_g1_3_17244;
  assign net_17245 = seg_3_18_local_g1_4_17245;
  assign net_17246 = seg_3_18_local_g1_5_17246;
  assign net_17248 = seg_3_18_local_g1_7_17248;
  assign net_17249 = seg_3_18_local_g2_0_17249;
  assign net_17253 = seg_3_18_local_g2_4_17253;
  assign net_17259 = seg_3_18_local_g3_2_17259;
  assign net_17364 = seg_3_19_local_g1_0_17364;
  assign net_17373 = seg_3_19_local_g2_1_17373;
  assign net_17504 = seg_3_20_local_g3_1_17504;
  assign net_17613 = seg_3_21_local_g1_3_17613;
  assign net_17620 = seg_3_21_local_g2_2_17620;
  assign net_17745 = seg_3_22_local_g2_4_17745;
  assign net_18935 = seg_4_1_local_g0_2_18935;
  assign net_18936 = seg_4_1_local_g0_3_18936;
  assign net_18940 = seg_4_1_local_g0_7_18940;
  assign net_18942 = seg_4_1_local_g1_1_18942;
  assign net_18943 = seg_4_1_local_g1_2_18943;
  assign net_18944 = seg_4_1_local_g1_3_18944;
  assign net_18945 = seg_4_1_local_g1_4_18945;
  assign net_18946 = seg_4_1_local_g1_5_18946;
  assign net_18948 = seg_4_1_local_g1_7_18948;
  assign net_18949 = seg_4_1_local_g2_0_18949;
  assign net_18951 = seg_4_1_local_g2_2_18951;
  assign net_18952 = seg_4_1_local_g2_3_18952;
  assign net_18954 = seg_4_1_local_g2_5_18954;
  assign net_18960 = seg_4_1_local_g3_3_18960;
  assign net_18963 = seg_4_1_local_g3_6_18963;
  assign net_19098 = seg_4_2_local_g0_2_19098;
  assign net_19100 = seg_4_2_local_g0_4_19100;
  assign net_19102 = seg_4_2_local_g0_6_19102;
  assign net_19103 = seg_4_2_local_g0_7_19103;
  assign net_19107 = seg_4_2_local_g1_3_19107;
  assign net_19108 = seg_4_2_local_g1_4_19108;
  assign net_19109 = seg_4_2_local_g1_5_19109;
  assign net_19110 = seg_4_2_local_g1_6_19110;
  assign net_19113 = seg_4_2_local_g2_1_19113;
  assign net_19114 = seg_4_2_local_g2_2_19114;
  assign net_19117 = seg_4_2_local_g2_5_19117;
  assign net_19118 = seg_4_2_local_g2_6_19118;
  assign net_19119 = seg_4_2_local_g2_7_19119;
  assign net_19122 = seg_4_2_local_g3_2_19122;
  assign net_19123 = seg_4_2_local_g3_3_19123;
  assign net_19124 = seg_4_2_local_g3_4_19124;
  assign net_19126 = seg_4_2_local_g3_6_19126;
  assign net_19127 = seg_4_2_local_g3_7_19127;
  assign net_19219 = seg_4_3_local_g0_0_19219;
  assign net_19221 = seg_4_3_local_g0_2_19221;
  assign net_19222 = seg_4_3_local_g0_3_19222;
  assign net_19223 = seg_4_3_local_g0_4_19223;
  assign net_19224 = seg_4_3_local_g0_5_19224;
  assign net_19225 = seg_4_3_local_g0_6_19225;
  assign net_19230 = seg_4_3_local_g1_3_19230;
  assign net_19231 = seg_4_3_local_g1_4_19231;
  assign net_19232 = seg_4_3_local_g1_5_19232;
  assign net_19233 = seg_4_3_local_g1_6_19233;
  assign net_19234 = seg_4_3_local_g1_7_19234;
  assign net_19236 = seg_4_3_local_g2_1_19236;
  assign net_19237 = seg_4_3_local_g2_2_19237;
  assign net_19239 = seg_4_3_local_g2_4_19239;
  assign net_19240 = seg_4_3_local_g2_5_19240;
  assign net_19241 = seg_4_3_local_g2_6_19241;
  assign net_19242 = seg_4_3_local_g2_7_19242;
  assign net_19245 = seg_4_3_local_g3_2_19245;
  assign net_19247 = seg_4_3_local_g3_4_19247;
  assign net_19250 = seg_4_3_local_g3_7_19250;
  assign net_19346 = seg_4_4_local_g0_4_19346;
  assign net_19348 = seg_4_4_local_g0_6_19348;
  assign net_19350 = seg_4_4_local_g1_0_19350;
  assign net_19352 = seg_4_4_local_g1_2_19352;
  assign net_19353 = seg_4_4_local_g1_3_19353;
  assign net_19354 = seg_4_4_local_g1_4_19354;
  assign net_19356 = seg_4_4_local_g1_6_19356;
  assign net_19360 = seg_4_4_local_g2_2_19360;
  assign net_19361 = seg_4_4_local_g2_3_19361;
  assign net_19362 = seg_4_4_local_g2_4_19362;
  assign net_19365 = seg_4_4_local_g2_7_19365;
  assign net_19371 = seg_4_4_local_g3_5_19371;
  assign net_19373 = seg_4_4_local_g3_7_19373;
  assign net_19470 = seg_4_5_local_g0_5_19470;
  assign net_19471 = seg_4_5_local_g0_6_19471;
  assign net_19473 = seg_4_5_local_g1_0_19473;
  assign net_19474 = seg_4_5_local_g1_1_19474;
  assign net_19478 = seg_4_5_local_g1_5_19478;
  assign net_19479 = seg_4_5_local_g1_6_19479;
  assign net_19481 = seg_4_5_local_g2_0_19481;
  assign net_19483 = seg_4_5_local_g2_2_19483;
  assign net_19485 = seg_4_5_local_g2_4_19485;
  assign net_19488 = seg_4_5_local_g2_7_19488;
  assign net_19492 = seg_4_5_local_g3_3_19492;
  assign net_19493 = seg_4_5_local_g3_4_19493;
  assign net_19494 = seg_4_5_local_g3_5_19494;
  assign net_19495 = seg_4_5_local_g3_6_19495;
  assign net_19496 = seg_4_5_local_g3_7_19496;
  assign net_19588 = seg_4_6_local_g0_0_19588;
  assign net_19590 = seg_4_6_local_g0_2_19590;
  assign net_19591 = seg_4_6_local_g0_3_19591;
  assign net_19592 = seg_4_6_local_g0_4_19592;
  assign net_19595 = seg_4_6_local_g0_7_19595;
  assign net_19596 = seg_4_6_local_g1_0_19596;
  assign net_19599 = seg_4_6_local_g1_3_19599;
  assign net_19602 = seg_4_6_local_g1_6_19602;
  assign net_19603 = seg_4_6_local_g1_7_19603;
  assign net_19604 = seg_4_6_local_g2_0_19604;
  assign net_19612 = seg_4_6_local_g3_0_19612;
  assign net_19615 = seg_4_6_local_g3_3_19615;
  assign net_19712 = seg_4_7_local_g0_1_19712;
  assign net_19715 = seg_4_7_local_g0_4_19715;
  assign net_19718 = seg_4_7_local_g0_7_19718;
  assign net_19720 = seg_4_7_local_g1_1_19720;
  assign net_19721 = seg_4_7_local_g1_2_19721;
  assign net_19724 = seg_4_7_local_g1_5_19724;
  assign net_19725 = seg_4_7_local_g1_6_19725;
  assign net_19726 = seg_4_7_local_g1_7_19726;
  assign net_19729 = seg_4_7_local_g2_2_19729;
  assign net_19731 = seg_4_7_local_g2_4_19731;
  assign net_19732 = seg_4_7_local_g2_5_19732;
  assign net_19734 = seg_4_7_local_g2_7_19734;
  assign net_19735 = seg_4_7_local_g3_0_19735;
  assign net_19736 = seg_4_7_local_g3_1_19736;
  assign net_19737 = seg_4_7_local_g3_2_19737;
  assign net_19738 = seg_4_7_local_g3_3_19738;
  assign net_19740 = seg_4_7_local_g3_5_19740;
  assign net_19742 = seg_4_7_local_g3_7_19742;
  assign net_19838 = seg_4_8_local_g0_4_19838;
  assign net_19848 = seg_4_8_local_g1_6_19848;
  assign net_19852 = seg_4_8_local_g2_2_19852;
  assign net_19854 = seg_4_8_local_g2_4_19854;
  assign net_19856 = seg_4_8_local_g2_6_19856;
  assign net_19859 = seg_4_8_local_g3_1_19859;
  assign net_19861 = seg_4_8_local_g3_3_19861;
  assign net_19863 = seg_4_8_local_g3_5_19863;
  assign net_19865 = seg_4_8_local_g3_7_19865;
  assign net_19960 = seg_4_9_local_g0_3_19960;
  assign net_19972 = seg_4_9_local_g1_7_19972;
  assign net_20101 = seg_4_10_local_g2_5_20101;
  assign net_20111 = seg_4_10_local_g3_7_20111;
  assign net_20204 = seg_4_11_local_g0_1_20204;
  assign net_20205 = seg_4_11_local_g0_2_20205;
  assign net_20207 = seg_4_11_local_g0_4_20207;
  assign net_20213 = seg_4_11_local_g1_2_20213;
  assign net_20215 = seg_4_11_local_g1_4_20215;
  assign net_20220 = seg_4_11_local_g2_1_20220;
  assign net_20228 = seg_4_11_local_g3_1_20228;
  assign net_20232 = seg_4_11_local_g3_5_20232;
  assign net_20333 = seg_4_12_local_g0_7_20333;
  assign net_20337 = seg_4_12_local_g1_3_20337;
  assign net_20341 = seg_4_12_local_g1_7_20341;
  assign net_20344 = seg_4_12_local_g2_2_20344;
  assign net_20348 = seg_4_12_local_g2_6_20348;
  assign net_20350 = seg_4_12_local_g3_0_20350;
  assign net_20352 = seg_4_12_local_g3_2_20352;
  assign net_20449 = seg_4_13_local_g0_0_20449;
  assign net_20450 = seg_4_13_local_g0_1_20450;
  assign net_20452 = seg_4_13_local_g0_3_20452;
  assign net_20453 = seg_4_13_local_g0_4_20453;
  assign net_20455 = seg_4_13_local_g0_6_20455;
  assign net_20459 = seg_4_13_local_g1_2_20459;
  assign net_20460 = seg_4_13_local_g1_3_20460;
  assign net_20466 = seg_4_13_local_g2_1_20466;
  assign net_20470 = seg_4_13_local_g2_5_20470;
  assign net_20471 = seg_4_13_local_g2_6_20471;
  assign net_20472 = seg_4_13_local_g2_7_20472;
  assign net_20476 = seg_4_13_local_g3_3_20476;
  assign net_20477 = seg_4_13_local_g3_4_20477;
  assign net_20478 = seg_4_13_local_g3_5_20478;
  assign net_20584 = seg_4_14_local_g1_4_20584;
  assign net_20591 = seg_4_14_local_g2_3_20591;
  assign net_20593 = seg_4_14_local_g2_5_20593;
  assign net_20596 = seg_4_14_local_g3_0_20596;
  assign net_20598 = seg_4_14_local_g3_2_20598;
  assign net_20601 = seg_4_14_local_g3_5_20601;
  assign net_20602 = seg_4_14_local_g3_6_20602;
  assign net_20695 = seg_4_15_local_g0_0_20695;
  assign net_20712 = seg_4_15_local_g2_1_20712;
  assign net_20713 = seg_4_15_local_g2_2_20713;
  assign net_20715 = seg_4_15_local_g2_4_20715;
  assign net_20717 = seg_4_15_local_g2_6_20717;
  assign net_20721 = seg_4_15_local_g3_2_20721;
  assign net_20725 = seg_4_15_local_g3_6_20725;
  assign net_20726 = seg_4_15_local_g3_7_20726;
  assign net_20818 = seg_4_16_local_g0_0_20818;
  assign net_20825 = seg_4_16_local_g0_7_20825;
  assign net_20831 = seg_4_16_local_g1_5_20831;
  assign net_20834 = seg_4_16_local_g2_0_20834;
  assign net_20841 = seg_4_16_local_g2_7_20841;
  assign net_20846 = seg_4_16_local_g3_4_20846;
  assign net_20942 = seg_4_17_local_g0_1_20942;
  assign net_20949 = seg_4_17_local_g1_0_20949;
  assign net_20952 = seg_4_17_local_g1_3_20952;
  assign net_20954 = seg_4_17_local_g1_5_20954;
  assign net_20955 = seg_4_17_local_g1_6_20955;
  assign net_20958 = seg_4_17_local_g2_1_20958;
  assign net_20967 = seg_4_17_local_g3_2_20967;
  assign net_21070 = seg_4_18_local_g0_6_21070;
  assign net_21075 = seg_4_18_local_g1_3_21075;
  assign net_21078 = seg_4_18_local_g1_6_21078;
  assign net_21088 = seg_4_18_local_g3_0_21088;
  assign net_21091 = seg_4_18_local_g3_3_21091;
  assign net_21192 = seg_4_19_local_g0_5_21192;
  assign net_21196 = seg_4_19_local_g1_1_21196;
  assign net_21205 = seg_4_19_local_g2_2_21205;
  assign net_21315 = seg_4_20_local_g0_5_21315;
  assign net_21317 = seg_4_20_local_g0_7_21317;
  assign net_21579 = seg_4_22_local_g2_7_21579;
  assign net_22721 = seg_5_0_local_g1_7_22721;
  assign net_22785 = seg_5_1_local_g2_5_22785;
  assign net_22790 = seg_5_1_local_g3_2_22790;
  assign net_22791 = seg_5_1_local_g3_3_22791;
  assign net_22944 = seg_5_2_local_g2_1_22944;
  assign net_22955 = seg_5_2_local_g3_4_22955;
  assign net_23055 = seg_5_3_local_g0_5_23055;
  assign net_23056 = seg_5_3_local_g0_6_23056;
  assign net_23061 = seg_5_3_local_g1_3_23061;
  assign net_23063 = seg_5_3_local_g1_5_23063;
  assign net_23069 = seg_5_3_local_g2_3_23069;
  assign net_23071 = seg_5_3_local_g2_5_23071;
  assign net_23077 = seg_5_3_local_g3_3_23077;
  assign net_23078 = seg_5_3_local_g3_4_23078;
  assign net_2315 = seg_0_11_local_g0_1_2315;
  assign net_23177 = seg_5_4_local_g0_4_23177;
  assign net_23179 = seg_5_4_local_g0_6_23179;
  assign net_23186 = seg_5_4_local_g1_5_23186;
  assign net_23188 = seg_5_4_local_g1_7_23188;
  assign net_23189 = seg_5_4_local_g2_0_23189;
  assign net_23190 = seg_5_4_local_g2_1_23190;
  assign net_23197 = seg_5_4_local_g3_0_23197;
  assign net_23198 = seg_5_4_local_g3_1_23198;
  assign net_23204 = seg_5_4_local_g3_7_23204;
  assign net_2322 = seg_0_11_local_g1_0_2322;
  assign net_2327 = seg_0_11_local_g1_5_2327;
  assign net_23299 = seg_5_5_local_g0_3_23299;
  assign net_2330 = seg_0_11_local_g2_0_2330;
  assign net_23301 = seg_5_5_local_g0_5_23301;
  assign net_23305 = seg_5_5_local_g1_1_23305;
  assign net_23306 = seg_5_5_local_g1_2_23306;
  assign net_23307 = seg_5_5_local_g1_3_23307;
  assign net_23308 = seg_5_5_local_g1_4_23308;
  assign net_2331 = seg_0_11_local_g2_1_2331;
  assign net_23310 = seg_5_5_local_g1_6_23310;
  assign net_2332 = seg_0_11_local_g2_2_2332;
  assign net_23327 = seg_5_5_local_g3_7_23327;
  assign net_2333 = seg_0_11_local_g2_3_2333;
  assign net_2334 = seg_0_11_local_g2_4_2334;
  assign net_2336 = seg_0_11_local_g2_6_2336;
  assign net_2337 = seg_0_11_local_g2_7_2337;
  assign net_2338 = seg_0_11_local_g3_0_2338;
  assign net_2339 = seg_0_11_local_g3_1_2339;
  assign net_2340 = seg_0_11_local_g3_2_2340;
  assign net_23419 = seg_5_6_local_g0_0_23419;
  assign net_2342 = seg_0_11_local_g3_4_2342;
  assign net_23421 = seg_5_6_local_g0_2_23421;
  assign net_23422 = seg_5_6_local_g0_3_23422;
  assign net_23423 = seg_5_6_local_g0_4_23423;
  assign net_23424 = seg_5_6_local_g0_5_23424;
  assign net_23425 = seg_5_6_local_g0_6_23425;
  assign net_23426 = seg_5_6_local_g0_7_23426;
  assign net_23427 = seg_5_6_local_g1_0_23427;
  assign net_2343 = seg_0_11_local_g3_5_2343;
  assign net_23436 = seg_5_6_local_g2_1_23436;
  assign net_23443 = seg_5_6_local_g3_0_23443;
  assign net_23445 = seg_5_6_local_g3_2_23445;
  assign net_23446 = seg_5_6_local_g3_3_23446;
  assign net_23448 = seg_5_6_local_g3_5_23448;
  assign net_2345 = seg_0_11_local_g3_7_2345;
  assign net_23547 = seg_5_7_local_g0_5_23547;
  assign net_23548 = seg_5_7_local_g0_6_23548;
  assign net_23551 = seg_5_7_local_g1_1_23551;
  assign net_23553 = seg_5_7_local_g1_3_23553;
  assign net_23554 = seg_5_7_local_g1_4_23554;
  assign net_23555 = seg_5_7_local_g1_5_23555;
  assign net_23556 = seg_5_7_local_g1_6_23556;
  assign net_23567 = seg_5_7_local_g3_1_23567;
  assign net_23571 = seg_5_7_local_g3_5_23571;
  assign net_23668 = seg_5_8_local_g0_3_23668;
  assign net_23670 = seg_5_8_local_g0_5_23670;
  assign net_23671 = seg_5_8_local_g0_6_23671;
  assign net_23672 = seg_5_8_local_g0_7_23672;
  assign net_23674 = seg_5_8_local_g1_1_23674;
  assign net_23676 = seg_5_8_local_g1_3_23676;
  assign net_23678 = seg_5_8_local_g1_5_23678;
  assign net_23682 = seg_5_8_local_g2_1_23682;
  assign net_23684 = seg_5_8_local_g2_3_23684;
  assign net_23687 = seg_5_8_local_g2_6_23687;
  assign net_23804 = seg_5_9_local_g2_0_23804;
  assign net_23805 = seg_5_9_local_g2_1_23805;
  assign net_23806 = seg_5_9_local_g2_2_23806;
  assign net_23807 = seg_5_9_local_g2_3_23807;
  assign net_23811 = seg_5_9_local_g2_7_23811;
  assign net_23812 = seg_5_9_local_g3_0_23812;
  assign net_23814 = seg_5_9_local_g3_2_23814;
  assign net_23817 = seg_5_9_local_g3_5_23817;
  assign net_23914 = seg_5_10_local_g0_3_23914;
  assign net_23916 = seg_5_10_local_g0_5_23916;
  assign net_23918 = seg_5_10_local_g0_7_23918;
  assign net_23920 = seg_5_10_local_g1_1_23920;
  assign net_23929 = seg_5_10_local_g2_2_23929;
  assign net_23933 = seg_5_10_local_g2_6_23933;
  assign net_23937 = seg_5_10_local_g3_2_23937;
  assign net_23939 = seg_5_10_local_g3_4_23939;
  assign net_24042 = seg_5_11_local_g1_0_24042;
  assign net_24049 = seg_5_11_local_g1_7_24049;
  assign net_24050 = seg_5_11_local_g2_0_24050;
  assign net_24052 = seg_5_11_local_g2_2_24052;
  assign net_24054 = seg_5_11_local_g2_4_24054;
  assign net_24058 = seg_5_11_local_g3_0_24058;
  assign net_24060 = seg_5_11_local_g3_2_24060;
  assign net_24062 = seg_5_11_local_g3_4_24062;
  assign net_24161 = seg_5_12_local_g0_4_24161;
  assign net_24164 = seg_5_12_local_g0_7_24164;
  assign net_24170 = seg_5_12_local_g1_5_24170;
  assign net_24173 = seg_5_12_local_g2_0_24173;
  assign net_24175 = seg_5_12_local_g2_2_24175;
  assign net_24177 = seg_5_12_local_g2_4_24177;
  assign net_24182 = seg_5_12_local_g3_1_24182;
  assign net_24184 = seg_5_12_local_g3_3_24184;
  assign net_24283 = seg_5_13_local_g0_3_24283;
  assign net_24286 = seg_5_13_local_g0_6_24286;
  assign net_24293 = seg_5_13_local_g1_5_24293;
  assign net_24296 = seg_5_13_local_g2_0_24296;
  assign net_24298 = seg_5_13_local_g2_2_24298;
  assign net_24300 = seg_5_13_local_g2_4_24300;
  assign net_24306 = seg_5_13_local_g3_2_24306;
  assign net_24310 = seg_5_13_local_g3_6_24310;
  assign net_24416 = seg_5_14_local_g1_5_24416;
  assign net_24421 = seg_5_14_local_g2_2_24421;
  assign net_24423 = seg_5_14_local_g2_4_24423;
  assign net_24428 = seg_5_14_local_g3_1_24428;
  assign net_24431 = seg_5_14_local_g3_4_24431;
  assign net_24432 = seg_5_14_local_g3_5_24432;
  assign net_24533 = seg_5_15_local_g0_7_24533;
  assign net_24535 = seg_5_15_local_g1_1_24535;
  assign net_24538 = seg_5_15_local_g1_4_24538;
  assign net_24548 = seg_5_15_local_g2_6_24548;
  assign net_24551 = seg_5_15_local_g3_1_24551;
  assign net_24553 = seg_5_15_local_g3_3_24553;
  assign net_24557 = seg_5_15_local_g3_7_24557;
  assign net_24649 = seg_5_16_local_g0_0_24649;
  assign net_24651 = seg_5_16_local_g0_2_24651;
  assign net_24653 = seg_5_16_local_g0_4_24653;
  assign net_24654 = seg_5_16_local_g0_5_24654;
  assign net_24656 = seg_5_16_local_g0_7_24656;
  assign net_24657 = seg_5_16_local_g1_0_24657;
  assign net_24658 = seg_5_16_local_g1_1_24658;
  assign net_24659 = seg_5_16_local_g1_2_24659;
  assign net_24660 = seg_5_16_local_g1_3_24660;
  assign net_24661 = seg_5_16_local_g1_4_24661;
  assign net_24662 = seg_5_16_local_g1_5_24662;
  assign net_24665 = seg_5_16_local_g2_0_24665;
  assign net_24675 = seg_5_16_local_g3_2_24675;
  assign net_24676 = seg_5_16_local_g3_3_24676;
  assign net_24680 = seg_5_16_local_g3_7_24680;
  assign net_24772 = seg_5_17_local_g0_0_24772;
  assign net_24773 = seg_5_17_local_g0_1_24773;
  assign net_24780 = seg_5_17_local_g1_0_24780;
  assign net_24783 = seg_5_17_local_g1_3_24783;
  assign net_24792 = seg_5_17_local_g2_4_24792;
  assign net_24895 = seg_5_18_local_g0_0_24895;
  assign net_24899 = seg_5_18_local_g0_4_24899;
  assign net_24925 = seg_5_18_local_g3_6_24925;
  assign net_25024 = seg_5_19_local_g0_6_25024;
  assign net_25038 = seg_5_19_local_g2_4_25038;
  assign net_2520 = seg_0_12_local_g0_0_2520;
  assign net_2521 = seg_0_12_local_g0_1_2521;
  assign net_2522 = seg_0_12_local_g0_2_2522;
  assign net_2523 = seg_0_12_local_g0_3_2523;
  assign net_2524 = seg_0_12_local_g0_4_2524;
  assign net_2526 = seg_0_12_local_g0_6_2526;
  assign net_2528 = seg_0_12_local_g1_0_2528;
  assign net_2529 = seg_0_12_local_g1_1_2529;
  assign net_2530 = seg_0_12_local_g1_2_2530;
  assign net_2531 = seg_0_12_local_g1_3_2531;
  assign net_2533 = seg_0_12_local_g1_5_2533;
  assign net_2534 = seg_0_12_local_g1_6_2534;
  assign net_2535 = seg_0_12_local_g1_7_2535;
  assign net_2544 = seg_0_12_local_g3_0_2544;
  assign net_2546 = seg_0_12_local_g3_2_2546;
  assign net_2548 = seg_0_12_local_g3_4_2548;
  assign net_26839 = seg_6_3_local_g0_2_26839;
  assign net_26841 = seg_6_3_local_g0_4_26841;
  assign net_26843 = seg_6_3_local_g0_6_26843;
  assign net_26844 = seg_6_3_local_g0_7_26844;
  assign net_26847 = seg_6_3_local_g1_2_26847;
  assign net_26849 = seg_6_3_local_g1_4_26849;
  assign net_26850 = seg_6_3_local_g1_5_26850;
  assign net_26853 = seg_6_3_local_g2_0_26853;
  assign net_26855 = seg_6_3_local_g2_2_26855;
  assign net_26856 = seg_6_3_local_g2_3_26856;
  assign net_26860 = seg_6_3_local_g2_7_26860;
  assign net_26861 = seg_6_3_local_g3_0_26861;
  assign net_26862 = seg_6_3_local_g3_1_26862;
  assign net_26866 = seg_6_3_local_g3_5_26866;
  assign net_26867 = seg_6_3_local_g3_6_26867;
  assign net_26939 = seg_6_4_local_g0_0_26939;
  assign net_26943 = seg_6_4_local_g0_4_26943;
  assign net_26944 = seg_6_4_local_g0_5_26944;
  assign net_26945 = seg_6_4_local_g0_6_26945;
  assign net_26949 = seg_6_4_local_g1_2_26949;
  assign net_26950 = seg_6_4_local_g1_3_26950;
  assign net_26951 = seg_6_4_local_g1_4_26951;
  assign net_26952 = seg_6_4_local_g1_5_26952;
  assign net_26955 = seg_6_4_local_g2_0_26955;
  assign net_26956 = seg_6_4_local_g2_1_26956;
  assign net_26957 = seg_6_4_local_g2_2_26957;
  assign net_26960 = seg_6_4_local_g2_5_26960;
  assign net_26961 = seg_6_4_local_g2_6_26961;
  assign net_26962 = seg_6_4_local_g2_7_26962;
  assign net_26964 = seg_6_4_local_g3_1_26964;
  assign net_26965 = seg_6_4_local_g3_2_26965;
  assign net_26968 = seg_6_4_local_g3_5_26968;
  assign net_26969 = seg_6_4_local_g3_6_26969;
  assign net_27467 = seg_6_9_local_g2_2_27467;
  assign net_27469 = seg_6_9_local_g2_4_27469;
  assign net_27471 = seg_6_9_local_g2_6_27471;
  assign net_27477 = seg_6_9_local_g3_4_27477;
  assign net_27569 = seg_6_10_local_g2_2_27569;
  assign net_27655 = seg_6_11_local_g0_2_27655;
  assign net_27657 = seg_6_11_local_g0_4_27657;
  assign net_27659 = seg_6_11_local_g0_6_27659;
  assign net_27665 = seg_6_11_local_g1_4_27665;
  assign net_27766 = seg_6_12_local_g1_3_27766;
  assign net_29752 = seg_7_0_local_g1_7_29752;
  assign net_29823 = seg_7_1_local_g3_4_29823;
  assign net_29961 = seg_7_2_local_g0_3_29961;
  assign net_29980 = seg_7_2_local_g2_6_29980;
  assign net_29983 = seg_7_2_local_g3_1_29983;
  assign net_30081 = seg_7_3_local_g0_0_30081;
  assign net_30091 = seg_7_3_local_g1_2_30091;
  assign net_30104 = seg_7_3_local_g2_7_30104;
  assign net_30112 = seg_7_3_local_g3_7_30112;
  assign net_30208 = seg_7_4_local_g0_4_30208;
  assign net_30211 = seg_7_4_local_g0_7_30211;
  assign net_30221 = seg_7_4_local_g2_1_30221;
  assign net_30224 = seg_7_4_local_g2_4_30224;
  assign net_30225 = seg_7_4_local_g2_5_30225;
  assign net_30232 = seg_7_4_local_g3_4_30232;
  assign net_30235 = seg_7_4_local_g3_7_30235;
  assign net_30329 = seg_7_5_local_g0_2_30329;
  assign net_30333 = seg_7_5_local_g0_6_30333;
  assign net_30336 = seg_7_5_local_g1_1_30336;
  assign net_30337 = seg_7_5_local_g1_2_30337;
  assign net_30341 = seg_7_5_local_g1_6_30341;
  assign net_30342 = seg_7_5_local_g1_7_30342;
  assign net_30343 = seg_7_5_local_g2_0_30343;
  assign net_30346 = seg_7_5_local_g2_3_30346;
  assign net_30348 = seg_7_5_local_g2_5_30348;
  assign net_30350 = seg_7_5_local_g2_7_30350;
  assign net_30354 = seg_7_5_local_g3_3_30354;
  assign net_30355 = seg_7_5_local_g3_4_30355;
  assign net_30358 = seg_7_5_local_g3_7_30358;
  assign net_30453 = seg_7_6_local_g0_3_30453;
  assign net_30455 = seg_7_6_local_g0_5_30455;
  assign net_30459 = seg_7_6_local_g1_1_30459;
  assign net_30460 = seg_7_6_local_g1_2_30460;
  assign net_30461 = seg_7_6_local_g1_3_30461;
  assign net_30463 = seg_7_6_local_g1_5_30463;
  assign net_30476 = seg_7_6_local_g3_2_30476;
  assign net_30477 = seg_7_6_local_g3_3_30477;
  assign net_30478 = seg_7_6_local_g3_4_30478;
  assign net_30481 = seg_7_6_local_g3_7_30481;
  assign net_30575 = seg_7_7_local_g0_2_30575;
  assign net_30576 = seg_7_7_local_g0_3_30576;
  assign net_30579 = seg_7_7_local_g0_6_30579;
  assign net_30580 = seg_7_7_local_g0_7_30580;
  assign net_30584 = seg_7_7_local_g1_3_30584;
  assign net_30591 = seg_7_7_local_g2_2_30591;
  assign net_30592 = seg_7_7_local_g2_3_30592;
  assign net_30601 = seg_7_7_local_g3_4_30601;
  assign net_30604 = seg_7_7_local_g3_7_30604;
  assign net_30696 = seg_7_8_local_g0_0_30696;
  assign net_30702 = seg_7_8_local_g0_6_30702;
  assign net_30704 = seg_7_8_local_g1_0_30704;
  assign net_30712 = seg_7_8_local_g2_0_30712;
  assign net_30718 = seg_7_8_local_g2_6_30718;
  assign net_30720 = seg_7_8_local_g3_0_30720;
  assign net_30724 = seg_7_8_local_g3_4_30724;
  assign net_30726 = seg_7_8_local_g3_6_30726;
  assign net_30820 = seg_7_9_local_g0_1_30820;
  assign net_30828 = seg_7_9_local_g1_1_30828;
  assign net_30830 = seg_7_9_local_g1_3_30830;
  assign net_30831 = seg_7_9_local_g1_4_30831;
  assign net_30836 = seg_7_9_local_g2_1_30836;
  assign net_30841 = seg_7_9_local_g2_6_30841;
  assign net_30848 = seg_7_9_local_g3_5_30848;
  assign net_30946 = seg_7_10_local_g0_4_30946;
  assign net_30950 = seg_7_10_local_g1_0_30950;
  assign net_30958 = seg_7_10_local_g2_0_30958;
  assign net_30959 = seg_7_10_local_g2_1_30959;
  assign net_30963 = seg_7_10_local_g2_5_30963;
  assign net_30967 = seg_7_10_local_g3_1_30967;
  assign net_30969 = seg_7_10_local_g3_3_30969;
  assign net_31071 = seg_7_11_local_g0_6_31071;
  assign net_31076 = seg_7_11_local_g1_3_31076;
  assign net_31079 = seg_7_11_local_g1_6_31079;
  assign net_31084 = seg_7_11_local_g2_3_31084;
  assign net_31086 = seg_7_11_local_g2_5_31086;
  assign net_31087 = seg_7_11_local_g2_6_31087;
  assign net_31091 = seg_7_11_local_g3_2_31091;
  assign net_31095 = seg_7_11_local_g3_6_31095;
  assign net_31189 = seg_7_12_local_g0_1_31189;
  assign net_31190 = seg_7_12_local_g0_2_31190;
  assign net_31191 = seg_7_12_local_g0_3_31191;
  assign net_31192 = seg_7_12_local_g0_4_31192;
  assign net_31195 = seg_7_12_local_g0_7_31195;
  assign net_31196 = seg_7_12_local_g1_0_31196;
  assign net_31197 = seg_7_12_local_g1_1_31197;
  assign net_31198 = seg_7_12_local_g1_2_31198;
  assign net_31199 = seg_7_12_local_g1_3_31199;
  assign net_31201 = seg_7_12_local_g1_5_31201;
  assign net_31203 = seg_7_12_local_g1_7_31203;
  assign net_31207 = seg_7_12_local_g2_3_31207;
  assign net_31214 = seg_7_12_local_g3_2_31214;
  assign net_31217 = seg_7_12_local_g3_5_31217;
  assign net_31312 = seg_7_13_local_g0_1_31312;
  assign net_31313 = seg_7_13_local_g0_2_31313;
  assign net_31314 = seg_7_13_local_g0_3_31314;
  assign net_31315 = seg_7_13_local_g0_4_31315;
  assign net_31319 = seg_7_13_local_g1_0_31319;
  assign net_31322 = seg_7_13_local_g1_3_31322;
  assign net_31331 = seg_7_13_local_g2_4_31331;
  assign net_31340 = seg_7_13_local_g3_5_31340;
  assign net_31444 = seg_7_14_local_g1_2_31444;
  assign net_31445 = seg_7_14_local_g1_3_31445;
  assign net_31448 = seg_7_14_local_g1_6_31448;
  assign net_31459 = seg_7_14_local_g3_1_31459;
  assign net_31557 = seg_7_15_local_g0_0_31557;
  assign net_31558 = seg_7_15_local_g0_1_31558;
  assign net_31559 = seg_7_15_local_g0_2_31559;
  assign net_31561 = seg_7_15_local_g0_4_31561;
  assign net_31562 = seg_7_15_local_g0_5_31562;
  assign net_31563 = seg_7_15_local_g0_6_31563;
  assign net_31564 = seg_7_15_local_g0_7_31564;
  assign net_31565 = seg_7_15_local_g1_0_31565;
  assign net_31566 = seg_7_15_local_g1_1_31566;
  assign net_31567 = seg_7_15_local_g1_2_31567;
  assign net_31568 = seg_7_15_local_g1_3_31568;
  assign net_31569 = seg_7_15_local_g1_4_31569;
  assign net_31570 = seg_7_15_local_g1_5_31570;
  assign net_31571 = seg_7_15_local_g1_6_31571;
  assign net_31572 = seg_7_15_local_g1_7_31572;
  assign net_31573 = seg_7_15_local_g2_0_31573;
  assign net_31574 = seg_7_15_local_g2_1_31574;
  assign net_31575 = seg_7_15_local_g2_2_31575;
  assign net_31577 = seg_7_15_local_g2_4_31577;
  assign net_31578 = seg_7_15_local_g2_5_31578;
  assign net_31582 = seg_7_15_local_g3_1_31582;
  assign net_31583 = seg_7_15_local_g3_2_31583;
  assign net_31584 = seg_7_15_local_g3_3_31584;
  assign net_31585 = seg_7_15_local_g3_4_31585;
  assign net_31586 = seg_7_15_local_g3_5_31586;
  assign net_31696 = seg_7_16_local_g2_0_31696;
  assign net_31699 = seg_7_16_local_g2_3_31699;
  assign net_31701 = seg_7_16_local_g2_5_31701;
  assign net_31709 = seg_7_16_local_g3_5_31709;
  assign net_31711 = seg_7_16_local_g3_7_31711;
  assign net_31805 = seg_7_17_local_g0_2_31805;
  assign net_31806 = seg_7_17_local_g0_3_31806;
  assign net_31807 = seg_7_17_local_g0_4_31807;
  assign net_31808 = seg_7_17_local_g0_5_31808;
  assign net_31811 = seg_7_17_local_g1_0_31811;
  assign net_31812 = seg_7_17_local_g1_1_31812;
  assign net_31813 = seg_7_17_local_g1_2_31813;
  assign net_31814 = seg_7_17_local_g1_3_31814;
  assign net_31816 = seg_7_17_local_g1_5_31816;
  assign net_31817 = seg_7_17_local_g1_6_31817;
  assign net_31818 = seg_7_17_local_g1_7_31818;
  assign net_31824 = seg_7_17_local_g2_5_31824;
  assign net_31832 = seg_7_17_local_g3_5_31832;
  assign net_31833 = seg_7_17_local_g3_6_31833;
  assign net_31932 = seg_7_18_local_g0_6_31932;
  assign net_31934 = seg_7_18_local_g1_0_31934;
  assign net_31937 = seg_7_18_local_g1_3_31937;
  assign net_31939 = seg_7_18_local_g1_5_31939;
  assign net_31954 = seg_7_18_local_g3_4_31954;
  assign net_31956 = seg_7_18_local_g3_6_31956;
  assign net_32065 = seg_7_19_local_g2_0_32065;
  assign net_32070 = seg_7_19_local_g2_5_32070;
  assign net_32072 = seg_7_19_local_g2_7_32072;
  assign net_32074 = seg_7_19_local_g3_1_32074;
  assign net_33572 = seg_8_0_local_g0_4_33572;
  assign net_33635 = seg_8_1_local_g1_1_33635;
  assign net_33644 = seg_8_1_local_g2_2_33644;
  assign net_33646 = seg_8_1_local_g2_4_33646;
  assign net_33648 = seg_8_1_local_g2_6_33648;
  assign net_33652 = seg_8_1_local_g3_2_33652;
  assign net_3380 = seg_0_16_local_g0_6_3380;
  assign net_33812 = seg_8_2_local_g2_7_33812;
  assign net_33813 = seg_8_2_local_g3_0_33813;
  assign net_33818 = seg_8_2_local_g3_5_33818;
  assign net_3382 = seg_0_16_local_g1_0_3382;
  assign net_3383 = seg_0_16_local_g1_1_3383;
  assign net_3385 = seg_0_16_local_g1_3_3385;
  assign net_3386 = seg_0_16_local_g1_4_3386;
  assign net_3388 = seg_0_16_local_g1_6_3388;
  assign net_3389 = seg_0_16_local_g1_7_3389;
  assign net_3390 = seg_0_16_local_g2_0_3390;
  assign net_33914 = seg_8_3_local_g0_2_33914;
  assign net_33917 = seg_8_3_local_g0_5_33917;
  assign net_33918 = seg_8_3_local_g0_6_33918;
  assign net_3392 = seg_0_16_local_g2_2_3392;
  assign net_3393 = seg_0_16_local_g2_3_3393;
  assign net_33931 = seg_8_3_local_g2_3_33931;
  assign net_33933 = seg_8_3_local_g2_5_33933;
  assign net_33934 = seg_8_3_local_g2_6_33934;
  assign net_33935 = seg_8_3_local_g2_7_33935;
  assign net_33937 = seg_8_3_local_g3_1_33937;
  assign net_3394 = seg_0_16_local_g2_4_3394;
  assign net_33941 = seg_8_3_local_g3_5_33941;
  assign net_3395 = seg_0_16_local_g2_5_3395;
  assign net_3397 = seg_0_16_local_g2_7_3397;
  assign net_3399 = seg_0_16_local_g3_1_3399;
  assign net_3400 = seg_0_16_local_g3_2_3400;
  assign net_3402 = seg_0_16_local_g3_4_3402;
  assign net_34038 = seg_8_4_local_g0_3_34038;
  assign net_34040 = seg_8_4_local_g0_5_34040;
  assign net_34045 = seg_8_4_local_g1_2_34045;
  assign net_34053 = seg_8_4_local_g2_2_34053;
  assign net_34055 = seg_8_4_local_g2_4_34055;
  assign net_34056 = seg_8_4_local_g2_5_34056;
  assign net_34064 = seg_8_4_local_g3_5_34064;
  assign net_34160 = seg_8_5_local_g0_2_34160;
  assign net_34167 = seg_8_5_local_g1_1_34167;
  assign net_34171 = seg_8_5_local_g1_5_34171;
  assign net_34179 = seg_8_5_local_g2_5_34179;
  assign net_34181 = seg_8_5_local_g2_7_34181;
  assign net_34185 = seg_8_5_local_g3_3_34185;
  assign net_34186 = seg_8_5_local_g3_4_34186;
  assign net_34187 = seg_8_5_local_g3_5_34187;
  assign net_34189 = seg_8_5_local_g3_7_34189;
  assign net_34284 = seg_8_6_local_g0_3_34284;
  assign net_34286 = seg_8_6_local_g0_5_34286;
  assign net_34294 = seg_8_6_local_g1_5_34294;
  assign net_34298 = seg_8_6_local_g2_1_34298;
  assign net_34300 = seg_8_6_local_g2_3_34300;
  assign net_34304 = seg_8_6_local_g2_7_34304;
  assign net_34306 = seg_8_6_local_g3_1_34306;
  assign net_34406 = seg_8_7_local_g0_2_34406;
  assign net_34409 = seg_8_7_local_g0_5_34409;
  assign net_34418 = seg_8_7_local_g1_6_34418;
  assign net_34528 = seg_8_8_local_g0_1_34528;
  assign net_34529 = seg_8_8_local_g0_2_34529;
  assign net_34531 = seg_8_8_local_g0_4_34531;
  assign net_34532 = seg_8_8_local_g0_5_34532;
  assign net_34534 = seg_8_8_local_g0_7_34534;
  assign net_34539 = seg_8_8_local_g1_4_34539;
  assign net_34540 = seg_8_8_local_g1_5_34540;
  assign net_34541 = seg_8_8_local_g1_6_34541;
  assign net_34542 = seg_8_8_local_g1_7_34542;
  assign net_34544 = seg_8_8_local_g2_1_34544;
  assign net_34547 = seg_8_8_local_g2_4_34547;
  assign net_34552 = seg_8_8_local_g3_1_34552;
  assign net_34553 = seg_8_8_local_g3_2_34553;
  assign net_34558 = seg_8_8_local_g3_7_34558;
  assign net_34652 = seg_8_9_local_g0_2_34652;
  assign net_34662 = seg_8_9_local_g1_4_34662;
  assign net_34664 = seg_8_9_local_g1_6_34664;
  assign net_34665 = seg_8_9_local_g1_7_34665;
  assign net_34668 = seg_8_9_local_g2_2_34668;
  assign net_34672 = seg_8_9_local_g2_6_34672;
  assign net_34676 = seg_8_9_local_g3_2_34676;
  assign net_34678 = seg_8_9_local_g3_4_34678;
  assign net_34773 = seg_8_10_local_g0_0_34773;
  assign net_34788 = seg_8_10_local_g1_7_34788;
  assign net_34791 = seg_8_10_local_g2_2_34791;
  assign net_34904 = seg_8_11_local_g1_0_34904;
  assign net_34906 = seg_8_11_local_g1_2_34906;
  assign net_34908 = seg_8_11_local_g1_4_34908;
  assign net_34916 = seg_8_11_local_g2_4_34916;
  assign net_34918 = seg_8_11_local_g2_6_34918;
  assign net_34920 = seg_8_11_local_g3_0_34920;
  assign net_34922 = seg_8_11_local_g3_2_34922;
  assign net_34926 = seg_8_11_local_g3_6_34926;
  assign net_35021 = seg_8_12_local_g0_2_35021;
  assign net_35023 = seg_8_12_local_g0_4_35023;
  assign net_35028 = seg_8_12_local_g1_1_35028;
  assign net_35030 = seg_8_12_local_g1_3_35030;
  assign net_35032 = seg_8_12_local_g1_5_35032;
  assign net_35033 = seg_8_12_local_g1_6_35033;
  assign net_35034 = seg_8_12_local_g1_7_35034;
  assign net_35035 = seg_8_12_local_g2_0_35035;
  assign net_35040 = seg_8_12_local_g2_5_35040;
  assign net_35154 = seg_8_13_local_g1_4_35154;
  assign net_35158 = seg_8_13_local_g2_0_35158;
  assign net_35161 = seg_8_13_local_g2_3_35161;
  assign net_35168 = seg_8_13_local_g3_2_35168;
  assign net_35170 = seg_8_13_local_g3_4_35170;
  assign net_35172 = seg_8_13_local_g3_6_35172;
  assign net_35173 = seg_8_13_local_g3_7_35173;
  assign net_35269 = seg_8_14_local_g0_4_35269;
  assign net_35273 = seg_8_14_local_g1_0_35273;
  assign net_35276 = seg_8_14_local_g1_3_35276;
  assign net_35281 = seg_8_14_local_g2_0_35281;
  assign net_35282 = seg_8_14_local_g2_1_35282;
  assign net_35388 = seg_8_15_local_g0_0_35388;
  assign net_35390 = seg_8_15_local_g0_2_35390;
  assign net_35391 = seg_8_15_local_g0_3_35391;
  assign net_35392 = seg_8_15_local_g0_4_35392;
  assign net_35394 = seg_8_15_local_g0_6_35394;
  assign net_35396 = seg_8_15_local_g1_0_35396;
  assign net_35397 = seg_8_15_local_g1_1_35397;
  assign net_35399 = seg_8_15_local_g1_3_35399;
  assign net_35400 = seg_8_15_local_g1_4_35400;
  assign net_35401 = seg_8_15_local_g1_5_35401;
  assign net_35402 = seg_8_15_local_g1_6_35402;
  assign net_35403 = seg_8_15_local_g1_7_35403;
  assign net_35404 = seg_8_15_local_g2_0_35404;
  assign net_35405 = seg_8_15_local_g2_1_35405;
  assign net_35406 = seg_8_15_local_g2_2_35406;
  assign net_35407 = seg_8_15_local_g2_3_35407;
  assign net_35410 = seg_8_15_local_g2_6_35410;
  assign net_35413 = seg_8_15_local_g3_1_35413;
  assign net_35414 = seg_8_15_local_g3_2_35414;
  assign net_35415 = seg_8_15_local_g3_3_35415;
  assign net_35416 = seg_8_15_local_g3_4_35416;
  assign net_35417 = seg_8_15_local_g3_5_35417;
  assign net_35419 = seg_8_15_local_g3_7_35419;
  assign net_35513 = seg_8_16_local_g0_2_35513;
  assign net_35515 = seg_8_16_local_g0_4_35515;
  assign net_35519 = seg_8_16_local_g1_0_35519;
  assign net_35522 = seg_8_16_local_g1_3_35522;
  assign net_35524 = seg_8_16_local_g1_5_35524;
  assign net_35525 = seg_8_16_local_g1_6_35525;
  assign net_35526 = seg_8_16_local_g1_7_35526;
  assign net_35528 = seg_8_16_local_g2_1_35528;
  assign net_35530 = seg_8_16_local_g2_3_35530;
  assign net_35533 = seg_8_16_local_g2_6_35533;
  assign net_35535 = seg_8_16_local_g3_0_35535;
  assign net_35536 = seg_8_16_local_g3_1_35536;
  assign net_3580 = seg_0_17_local_g0_0_3580;
  assign net_3582 = seg_0_17_local_g0_2_3582;
  assign net_3583 = seg_0_17_local_g0_3_3583;
  assign net_3585 = seg_0_17_local_g0_5_3585;
  assign net_3587 = seg_0_17_local_g0_7_3587;
  assign net_3589 = seg_0_17_local_g1_1_3589;
  assign net_3590 = seg_0_17_local_g1_2_3590;
  assign net_3592 = seg_0_17_local_g1_4_3592;
  assign net_3594 = seg_0_17_local_g1_6_3594;
  assign net_3595 = seg_0_17_local_g1_7_3595;
  assign net_3597 = seg_0_17_local_g2_1_3597;
  assign net_3598 = seg_0_17_local_g2_2_3598;
  assign net_3600 = seg_0_17_local_g2_4_3600;
  assign net_3606 = seg_0_17_local_g3_2_3606;
  assign net_3607 = seg_0_17_local_g3_3_3607;
  assign net_3611 = seg_0_17_local_g3_7_3611;
  assign net_37403 = seg_9_0_local_g0_4_37403;
  assign net_37406 = seg_9_0_local_g0_7_37406;
  assign net_37457 = seg_9_1_local_g0_0_37457;
  assign net_37462 = seg_9_1_local_g0_5_37462;
  assign net_37464 = seg_9_1_local_g0_7_37464;
  assign net_37468 = seg_9_1_local_g1_3_37468;
  assign net_37480 = seg_9_1_local_g2_7_37480;
  assign net_37631 = seg_9_2_local_g1_3_37631;
  assign net_37633 = seg_9_2_local_g1_5_37633;
  assign net_37743 = seg_9_3_local_g0_0_37743;
  assign net_37746 = seg_9_3_local_g0_3_37746;
  assign net_37749 = seg_9_3_local_g0_6_37749;
  assign net_37752 = seg_9_3_local_g1_1_37752;
  assign net_37754 = seg_9_3_local_g1_3_37754;
  assign net_37762 = seg_9_3_local_g2_3_37762;
  assign net_37868 = seg_9_4_local_g0_2_37868;
  assign net_37870 = seg_9_4_local_g0_4_37870;
  assign net_37872 = seg_9_4_local_g0_6_37872;
  assign net_37873 = seg_9_4_local_g0_7_37873;
  assign net_37876 = seg_9_4_local_g1_2_37876;
  assign net_37880 = seg_9_4_local_g1_6_37880;
  assign net_37884 = seg_9_4_local_g2_2_37884;
  assign net_37885 = seg_9_4_local_g2_3_37885;
  assign net_37895 = seg_9_4_local_g3_5_37895;
  assign net_37989 = seg_9_5_local_g0_0_37989;
  assign net_37995 = seg_9_5_local_g0_6_37995;
  assign net_37997 = seg_9_5_local_g1_0_37997;
  assign net_37998 = seg_9_5_local_g1_1_37998;
  assign net_38008 = seg_9_5_local_g2_3_38008;
  assign net_38011 = seg_9_5_local_g2_6_38011;
  assign net_38016 = seg_9_5_local_g3_3_38016;
  assign net_38118 = seg_9_6_local_g0_6_38118;
  assign net_38119 = seg_9_6_local_g0_7_38119;
  assign net_38120 = seg_9_6_local_g1_0_38120;
  assign net_38127 = seg_9_6_local_g1_7_38127;
  assign net_38236 = seg_9_7_local_g0_1_38236;
  assign net_38240 = seg_9_7_local_g0_5_38240;
  assign net_38242 = seg_9_7_local_g0_7_38242;
  assign net_38244 = seg_9_7_local_g1_1_38244;
  assign net_38246 = seg_9_7_local_g1_3_38246;
  assign net_38249 = seg_9_7_local_g1_6_38249;
  assign net_38253 = seg_9_7_local_g2_2_38253;
  assign net_38255 = seg_9_7_local_g2_4_38255;
  assign net_38256 = seg_9_7_local_g2_5_38256;
  assign net_38359 = seg_9_8_local_g0_1_38359;
  assign net_38361 = seg_9_8_local_g0_3_38361;
  assign net_38363 = seg_9_8_local_g0_5_38363;
  assign net_38364 = seg_9_8_local_g0_6_38364;
  assign net_38365 = seg_9_8_local_g0_7_38365;
  assign net_38368 = seg_9_8_local_g1_2_38368;
  assign net_38370 = seg_9_8_local_g1_4_38370;
  assign net_38373 = seg_9_8_local_g1_7_38373;
  assign net_38375 = seg_9_8_local_g2_1_38375;
  assign net_38380 = seg_9_8_local_g2_6_38380;
  assign net_38484 = seg_9_9_local_g0_3_38484;
  assign net_38485 = seg_9_9_local_g0_4_38485;
  assign net_38486 = seg_9_9_local_g0_5_38486;
  assign net_38487 = seg_9_9_local_g0_6_38487;
  assign net_38491 = seg_9_9_local_g1_2_38491;
  assign net_38494 = seg_9_9_local_g1_5_38494;
  assign net_38495 = seg_9_9_local_g1_6_38495;
  assign net_38604 = seg_9_10_local_g0_0_38604;
  assign net_38608 = seg_9_10_local_g0_4_38608;
  assign net_38614 = seg_9_10_local_g1_2_38614;
  assign net_38615 = seg_9_10_local_g1_3_38615;
  assign net_38616 = seg_9_10_local_g1_4_38616;
  assign net_38624 = seg_9_10_local_g2_4_38624;
  assign net_38629 = seg_9_10_local_g3_1_38629;
  assign net_38632 = seg_9_10_local_g3_4_38632;
  assign net_38735 = seg_9_11_local_g1_0_38735;
  assign net_38738 = seg_9_11_local_g1_3_38738;
  assign net_38749 = seg_9_11_local_g2_6_38749;
  assign net_38852 = seg_9_12_local_g0_2_38852;
  assign net_38858 = seg_9_12_local_g1_0_38858;
  assign net_38873 = seg_9_12_local_g2_7_38873;
  assign net_38877 = seg_9_12_local_g3_3_38877;
  assign net_38879 = seg_9_12_local_g3_5_38879;
  assign net_38880 = seg_9_12_local_g3_6_38880;
  assign net_38982 = seg_9_13_local_g1_1_38982;
  assign net_38983 = seg_9_13_local_g1_2_38983;
  assign net_38984 = seg_9_13_local_g1_3_38984;
  assign net_38990 = seg_9_13_local_g2_1_38990;
  assign net_38991 = seg_9_13_local_g2_2_38991;
  assign net_39000 = seg_9_13_local_g3_3_39000;
  assign net_39003 = seg_9_13_local_g3_6_39003;
  assign net_39098 = seg_9_14_local_g0_2_39098;
  assign net_39099 = seg_9_14_local_g0_3_39099;
  assign net_39100 = seg_9_14_local_g0_4_39100;
  assign net_39107 = seg_9_14_local_g1_3_39107;
  assign net_39110 = seg_9_14_local_g1_6_39110;
  assign net_39114 = seg_9_14_local_g2_2_39114;
  assign net_39115 = seg_9_14_local_g2_3_39115;
  assign net_39118 = seg_9_14_local_g2_6_39118;
  assign net_39123 = seg_9_14_local_g3_3_39123;
  assign net_39126 = seg_9_14_local_g3_6_39126;
  assign net_39224 = seg_9_15_local_g0_5_39224;
  assign net_39228 = seg_9_15_local_g1_1_39228;
  assign net_39230 = seg_9_15_local_g1_3_39230;
  assign net_39231 = seg_9_15_local_g1_4_39231;
  assign net_39233 = seg_9_15_local_g1_6_39233;
  assign net_39234 = seg_9_15_local_g1_7_39234;
  assign net_39235 = seg_9_15_local_g2_0_39235;
  assign net_39236 = seg_9_15_local_g2_1_39236;
  assign net_39238 = seg_9_15_local_g2_3_39238;
  assign net_39244 = seg_9_15_local_g3_1_39244;
  assign net_39246 = seg_9_15_local_g3_3_39246;
  assign net_39247 = seg_9_15_local_g3_4_39247;
  assign net_39249 = seg_9_15_local_g3_6_39249;
  assign net_39344 = seg_9_16_local_g0_2_39344;
  assign net_39345 = seg_9_16_local_g0_3_39345;
  assign net_39348 = seg_9_16_local_g0_6_39348;
  assign net_39352 = seg_9_16_local_g1_2_39352;
  assign net_39360 = seg_9_16_local_g2_2_39360;
  assign net_39364 = seg_9_16_local_g2_6_39364;
  assign net_39466 = seg_9_17_local_g0_1_39466;
  assign net_39474 = seg_9_17_local_g1_1_39474;
  assign net_39476 = seg_9_17_local_g1_3_39476;
  assign net_39480 = seg_9_17_local_g1_7_39480;
  assign net_39481 = seg_9_17_local_g2_0_39481;
  assign net_39482 = seg_9_17_local_g2_1_39482;
  assign net_39483 = seg_9_17_local_g2_2_39483;
  assign net_39484 = seg_9_17_local_g2_3_39484;
  assign net_39492 = seg_9_17_local_g3_3_39492;
  assign net_39588 = seg_9_18_local_g0_0_39588;
  assign net_39589 = seg_9_18_local_g0_1_39589;
  assign net_39590 = seg_9_18_local_g0_2_39590;
  assign net_39591 = seg_9_18_local_g0_3_39591;
  assign net_39592 = seg_9_18_local_g0_4_39592;
  assign net_39594 = seg_9_18_local_g0_6_39594;
  assign net_39595 = seg_9_18_local_g0_7_39595;
  assign net_39596 = seg_9_18_local_g1_0_39596;
  assign net_39597 = seg_9_18_local_g1_1_39597;
  assign net_39598 = seg_9_18_local_g1_2_39598;
  assign net_39599 = seg_9_18_local_g1_3_39599;
  assign net_39600 = seg_9_18_local_g1_4_39600;
  assign net_39602 = seg_9_18_local_g1_6_39602;
  assign net_39603 = seg_9_18_local_g1_7_39603;
  assign net_39604 = seg_9_18_local_g2_0_39604;
  assign net_39608 = seg_9_18_local_g2_4_39608;
  assign net_39610 = seg_9_18_local_g2_6_39610;
  assign net_39612 = seg_9_18_local_g3_0_39612;
  assign net_39613 = seg_9_18_local_g3_1_39613;
  assign net_39615 = seg_9_18_local_g3_3_39615;
  assign net_39618 = seg_9_18_local_g3_6_39618;
  assign net_41289 = seg_10_1_local_g0_1_41289;
  assign net_41292 = seg_10_1_local_g0_4_41292;
  assign net_41293 = seg_10_1_local_g0_5_41293;
  assign net_41294 = seg_10_1_local_g0_6_41294;
  assign net_41299 = seg_10_1_local_g1_3_41299;
  assign net_41302 = seg_10_1_local_g1_6_41302;
  assign net_41303 = seg_10_1_local_g1_7_41303;
  assign net_41309 = seg_10_1_local_g2_5_41309;
  assign net_41452 = seg_10_2_local_g0_1_41452;
  assign net_41457 = seg_10_2_local_g0_6_41457;
  assign net_41458 = seg_10_2_local_g0_7_41458;
  assign net_41470 = seg_10_2_local_g2_3_41470;
  assign net_41474 = seg_10_2_local_g2_7_41474;
  assign net_41475 = seg_10_2_local_g3_0_41475;
  assign net_41477 = seg_10_2_local_g3_2_41477;
  assign net_41479 = seg_10_2_local_g3_4_41479;
  assign net_41584 = seg_10_3_local_g1_2_41584;
  assign net_41589 = seg_10_3_local_g1_7_41589;
  assign net_41593 = seg_10_3_local_g2_3_41593;
  assign net_41594 = seg_10_3_local_g2_4_41594;
  assign net_41595 = seg_10_3_local_g2_5_41595;
  assign net_41598 = seg_10_3_local_g3_0_41598;
  assign net_41603 = seg_10_3_local_g3_5_41603;
  assign net_41604 = seg_10_3_local_g3_6_41604;
  assign net_41703 = seg_10_4_local_g0_6_41703;
  assign net_41704 = seg_10_4_local_g0_7_41704;
  assign net_41706 = seg_10_4_local_g1_1_41706;
  assign net_41708 = seg_10_4_local_g1_3_41708;
  assign net_41710 = seg_10_4_local_g1_5_41710;
  assign net_41712 = seg_10_4_local_g1_7_41712;
  assign net_41714 = seg_10_4_local_g2_1_41714;
  assign net_41719 = seg_10_4_local_g2_6_41719;
  assign net_41724 = seg_10_4_local_g3_3_41724;
  assign net_41725 = seg_10_4_local_g3_4_41725;
  assign net_41727 = seg_10_4_local_g3_6_41727;
  assign net_41828 = seg_10_5_local_g1_0_41828;
  assign net_41832 = seg_10_5_local_g1_4_41832;
  assign net_41842 = seg_10_5_local_g2_6_41842;
  assign net_41846 = seg_10_5_local_g3_2_41846;
  assign net_41849 = seg_10_5_local_g3_5_41849;
  assign net_41953 = seg_10_6_local_g1_2_41953;
  assign net_41960 = seg_10_6_local_g2_1_41960;
  assign net_41968 = seg_10_6_local_g3_1_41968;
  assign net_42070 = seg_10_7_local_g0_4_42070;
  assign net_42072 = seg_10_7_local_g0_6_42072;
  assign net_42073 = seg_10_7_local_g0_7_42073;
  assign net_42074 = seg_10_7_local_g1_0_42074;
  assign net_42082 = seg_10_7_local_g2_0_42082;
  assign net_42091 = seg_10_7_local_g3_1_42091;
  assign net_42093 = seg_10_7_local_g3_3_42093;
  assign net_42193 = seg_10_8_local_g0_4_42193;
  assign net_42198 = seg_10_8_local_g1_1_42198;
  assign net_42199 = seg_10_8_local_g1_2_42199;
  assign net_42202 = seg_10_8_local_g1_5_42202;
  assign net_42203 = seg_10_8_local_g1_6_42203;
  assign net_42213 = seg_10_8_local_g3_0_42213;
  assign net_42218 = seg_10_8_local_g3_5_42218;
  assign net_42319 = seg_10_9_local_g0_7_42319;
  assign net_42436 = seg_10_10_local_g0_1_42436;
  assign net_42437 = seg_10_10_local_g0_2_42437;
  assign net_42439 = seg_10_10_local_g0_4_42439;
  assign net_42444 = seg_10_10_local_g1_1_42444;
  assign net_42445 = seg_10_10_local_g1_2_42445;
  assign net_42448 = seg_10_10_local_g1_5_42448;
  assign net_42454 = seg_10_10_local_g2_3_42454;
  assign net_42456 = seg_10_10_local_g2_5_42456;
  assign net_42558 = seg_10_11_local_g0_0_42558;
  assign net_42559 = seg_10_11_local_g0_1_42559;
  assign net_42560 = seg_10_11_local_g0_2_42560;
  assign net_42565 = seg_10_11_local_g0_7_42565;
  assign net_42567 = seg_10_11_local_g1_1_42567;
  assign net_42569 = seg_10_11_local_g1_3_42569;
  assign net_42572 = seg_10_11_local_g1_6_42572;
  assign net_42575 = seg_10_11_local_g2_1_42575;
  assign net_42576 = seg_10_11_local_g2_2_42576;
  assign net_42581 = seg_10_11_local_g2_7_42581;
  assign net_42588 = seg_10_11_local_g3_6_42588;
  assign net_42683 = seg_10_12_local_g0_2_42683;
  assign net_42692 = seg_10_12_local_g1_3_42692;
  assign net_42806 = seg_10_13_local_g0_2_42806;
  assign net_42810 = seg_10_13_local_g0_6_42810;
  assign net_42814 = seg_10_13_local_g1_2_42814;
  assign net_42927 = seg_10_14_local_g0_0_42927;
  assign net_42936 = seg_10_14_local_g1_1_42936;
  assign net_42951 = seg_10_14_local_g3_0_42951;
  assign net_42952 = seg_10_14_local_g3_1_42952;
  assign net_42953 = seg_10_14_local_g3_2_42953;
  assign net_42954 = seg_10_14_local_g3_3_42954;
  assign net_42955 = seg_10_14_local_g3_4_42955;
  assign net_43052 = seg_10_15_local_g0_2_43052;
  assign net_43053 = seg_10_15_local_g0_3_43053;
  assign net_43056 = seg_10_15_local_g0_6_43056;
  assign net_43061 = seg_10_15_local_g1_3_43061;
  assign net_43063 = seg_10_15_local_g1_5_43063;
  assign net_43065 = seg_10_15_local_g1_7_43065;
  assign net_43076 = seg_10_15_local_g3_2_43076;
  assign net_43077 = seg_10_15_local_g3_3_43077;
  assign net_43182 = seg_10_16_local_g1_1_43182;
  assign net_43187 = seg_10_16_local_g1_6_43187;
  assign net_43191 = seg_10_16_local_g2_2_43191;
  assign net_43192 = seg_10_16_local_g2_3_43192;
  assign net_43193 = seg_10_16_local_g2_4_43193;
  assign net_43196 = seg_10_16_local_g2_7_43196;
  assign net_43296 = seg_10_17_local_g0_0_43296;
  assign net_43298 = seg_10_17_local_g0_2_43298;
  assign net_43299 = seg_10_17_local_g0_3_43299;
  assign net_43300 = seg_10_17_local_g0_4_43300;
  assign net_43301 = seg_10_17_local_g0_5_43301;
  assign net_43302 = seg_10_17_local_g0_6_43302;
  assign net_43305 = seg_10_17_local_g1_1_43305;
  assign net_43307 = seg_10_17_local_g1_3_43307;
  assign net_43310 = seg_10_17_local_g1_6_43310;
  assign net_43315 = seg_10_17_local_g2_3_43315;
  assign net_43316 = seg_10_17_local_g2_4_43316;
  assign net_43319 = seg_10_17_local_g2_7_43319;
  assign net_43419 = seg_10_18_local_g0_0_43419;
  assign net_43421 = seg_10_18_local_g0_2_43421;
  assign net_43422 = seg_10_18_local_g0_3_43422;
  assign net_43425 = seg_10_18_local_g0_6_43425;
  assign net_43426 = seg_10_18_local_g0_7_43426;
  assign net_43428 = seg_10_18_local_g1_1_43428;
  assign net_43431 = seg_10_18_local_g1_4_43431;
  assign net_43432 = seg_10_18_local_g1_5_43432;
  assign net_43434 = seg_10_18_local_g1_7_43434;
  assign net_43435 = seg_10_18_local_g2_0_43435;
  assign net_43437 = seg_10_18_local_g2_2_43437;
  assign net_43438 = seg_10_18_local_g2_3_43438;
  assign net_43439 = seg_10_18_local_g2_4_43439;
  assign net_43441 = seg_10_18_local_g2_6_43441;
  assign net_43444 = seg_10_18_local_g3_1_43444;
  assign net_43448 = seg_10_18_local_g3_5_43448;
  assign net_43450 = seg_10_18_local_g3_7_43450;
  assign net_43544 = seg_10_19_local_g0_2_43544;
  assign net_43549 = seg_10_19_local_g0_7_43549;
  assign net_43551 = seg_10_19_local_g1_1_43551;
  assign net_43556 = seg_10_19_local_g1_6_43556;
  assign net_43557 = seg_10_19_local_g1_7_43557;
  assign net_43559 = seg_10_19_local_g2_1_43559;
  assign net_43568 = seg_10_19_local_g3_2_43568;
  assign net_43569 = seg_10_19_local_g3_3_43569;
  assign net_45135 = seg_11_1_local_g2_0_45135;
  assign net_45283 = seg_11_2_local_g0_1_45283;
  assign net_45296 = seg_11_2_local_g1_6_45296;
  assign net_45299 = seg_11_2_local_g2_1_45299;
  assign net_45300 = seg_11_2_local_g2_2_45300;
  assign net_45301 = seg_11_2_local_g2_3_45301;
  assign net_45304 = seg_11_2_local_g2_6_45304;
  assign net_45305 = seg_11_2_local_g2_7_45305;
  assign net_45308 = seg_11_2_local_g3_2_45308;
  assign net_45311 = seg_11_2_local_g3_5_45311;
  assign net_45312 = seg_11_2_local_g3_6_45312;
  assign net_45313 = seg_11_2_local_g3_7_45313;
  assign net_45408 = seg_11_3_local_g0_3_45408;
  assign net_45411 = seg_11_3_local_g0_6_45411;
  assign net_45412 = seg_11_3_local_g0_7_45412;
  assign net_45413 = seg_11_3_local_g1_0_45413;
  assign net_45414 = seg_11_3_local_g1_1_45414;
  assign net_45415 = seg_11_3_local_g1_2_45415;
  assign net_45417 = seg_11_3_local_g1_4_45417;
  assign net_45418 = seg_11_3_local_g1_5_45418;
  assign net_45420 = seg_11_3_local_g1_7_45420;
  assign net_45425 = seg_11_3_local_g2_4_45425;
  assign net_45427 = seg_11_3_local_g2_6_45427;
  assign net_45429 = seg_11_3_local_g3_0_45429;
  assign net_45430 = seg_11_3_local_g3_1_45430;
  assign net_45435 = seg_11_3_local_g3_6_45435;
  assign net_45529 = seg_11_4_local_g0_1_45529;
  assign net_45532 = seg_11_4_local_g0_4_45532;
  assign net_45533 = seg_11_4_local_g0_5_45533;
  assign net_45534 = seg_11_4_local_g0_6_45534;
  assign net_45538 = seg_11_4_local_g1_2_45538;
  assign net_45539 = seg_11_4_local_g1_3_45539;
  assign net_45541 = seg_11_4_local_g1_5_45541;
  assign net_45542 = seg_11_4_local_g1_6_45542;
  assign net_45543 = seg_11_4_local_g1_7_45543;
  assign net_45546 = seg_11_4_local_g2_2_45546;
  assign net_45554 = seg_11_4_local_g3_2_45554;
  assign net_45557 = seg_11_4_local_g3_5_45557;
  assign net_45653 = seg_11_5_local_g0_2_45653;
  assign net_45654 = seg_11_5_local_g0_3_45654;
  assign net_45658 = seg_11_5_local_g0_7_45658;
  assign net_45662 = seg_11_5_local_g1_3_45662;
  assign net_45663 = seg_11_5_local_g1_4_45663;
  assign net_45665 = seg_11_5_local_g1_6_45665;
  assign net_45666 = seg_11_5_local_g1_7_45666;
  assign net_45790 = seg_11_6_local_g2_0_45790;
  assign net_45791 = seg_11_6_local_g2_1_45791;
  assign net_45793 = seg_11_6_local_g2_3_45793;
  assign net_45796 = seg_11_6_local_g2_6_45796;
  assign net_45905 = seg_11_7_local_g1_0_45905;
  assign net_45909 = seg_11_7_local_g1_4_45909;
  assign net_45923 = seg_11_7_local_g3_2_45923;
  assign net_46021 = seg_11_8_local_g0_1_46021;
  assign net_46025 = seg_11_8_local_g0_5_46025;
  assign net_46028 = seg_11_8_local_g1_0_46028;
  assign net_46031 = seg_11_8_local_g1_3_46031;
  assign net_46033 = seg_11_8_local_g1_5_46033;
  assign net_46034 = seg_11_8_local_g1_6_46034;
  assign net_46040 = seg_11_8_local_g2_4_46040;
  assign net_46042 = seg_11_8_local_g2_6_46042;
  assign net_46043 = seg_11_8_local_g2_7_46043;
  assign net_46144 = seg_11_9_local_g0_1_46144;
  assign net_46154 = seg_11_9_local_g1_3_46154;
  assign net_46158 = seg_11_9_local_g1_7_46158;
  assign net_46268 = seg_11_10_local_g0_2_46268;
  assign net_46273 = seg_11_10_local_g0_7_46273;
  assign net_46283 = seg_11_10_local_g2_1_46283;
  assign net_46285 = seg_11_10_local_g2_3_46285;
  assign net_46389 = seg_11_11_local_g0_0_46389;
  assign net_46392 = seg_11_11_local_g0_3_46392;
  assign net_46395 = seg_11_11_local_g0_6_46395;
  assign net_46397 = seg_11_11_local_g1_0_46397;
  assign net_46401 = seg_11_11_local_g1_4_46401;
  assign net_46402 = seg_11_11_local_g1_5_46402;
  assign net_46403 = seg_11_11_local_g1_6_46403;
  assign net_46405 = seg_11_11_local_g2_0_46405;
  assign net_46409 = seg_11_11_local_g2_4_46409;
  assign net_46410 = seg_11_11_local_g2_5_46410;
  assign net_46414 = seg_11_11_local_g3_1_46414;
  assign net_46417 = seg_11_11_local_g3_4_46417;
  assign net_46512 = seg_11_12_local_g0_0_46512;
  assign net_46518 = seg_11_12_local_g0_6_46518;
  assign net_46519 = seg_11_12_local_g0_7_46519;
  assign net_46522 = seg_11_12_local_g1_2_46522;
  assign net_46523 = seg_11_12_local_g1_3_46523;
  assign net_46527 = seg_11_12_local_g1_7_46527;
  assign net_46529 = seg_11_12_local_g2_1_46529;
  assign net_46530 = seg_11_12_local_g2_2_46530;
  assign net_46535 = seg_11_12_local_g2_7_46535;
  assign net_46536 = seg_11_12_local_g3_0_46536;
  assign net_46538 = seg_11_12_local_g3_2_46538;
  assign net_46540 = seg_11_12_local_g3_4_46540;
  assign net_46543 = seg_11_12_local_g3_7_46543;
  assign net_46636 = seg_11_13_local_g0_1_46636;
  assign net_46644 = seg_11_13_local_g1_1_46644;
  assign net_46653 = seg_11_13_local_g2_2_46653;
  assign net_46655 = seg_11_13_local_g2_4_46655;
  assign net_46660 = seg_11_13_local_g3_1_46660;
  assign net_46661 = seg_11_13_local_g3_2_46661;
  assign net_46758 = seg_11_14_local_g0_0_46758;
  assign net_46761 = seg_11_14_local_g0_3_46761;
  assign net_46762 = seg_11_14_local_g0_4_46762;
  assign net_46768 = seg_11_14_local_g1_2_46768;
  assign net_46771 = seg_11_14_local_g1_5_46771;
  assign net_46785 = seg_11_14_local_g3_3_46785;
  assign net_46882 = seg_11_15_local_g0_1_46882;
  assign net_46885 = seg_11_15_local_g0_4_46885;
  assign net_46887 = seg_11_15_local_g0_6_46887;
  assign net_46896 = seg_11_15_local_g1_7_46896;
  assign net_46897 = seg_11_15_local_g2_0_46897;
  assign net_46899 = seg_11_15_local_g2_2_46899;
  assign net_46901 = seg_11_15_local_g2_4_46901;
  assign net_46902 = seg_11_15_local_g2_5_46902;
  assign net_46904 = seg_11_15_local_g2_7_46904;
  assign net_46910 = seg_11_15_local_g3_5_46910;
  assign net_46911 = seg_11_15_local_g3_6_46911;
  assign net_47008 = seg_11_16_local_g0_4_47008;
  assign net_47012 = seg_11_16_local_g1_0_47012;
  assign net_47013 = seg_11_16_local_g1_1_47013;
  assign net_47018 = seg_11_16_local_g1_6_47018;
  assign net_47022 = seg_11_16_local_g2_2_47022;
  assign net_47023 = seg_11_16_local_g2_3_47023;
  assign net_47030 = seg_11_16_local_g3_2_47030;
  assign net_47031 = seg_11_16_local_g3_3_47031;
  assign net_47033 = seg_11_16_local_g3_5_47033;
  assign net_47128 = seg_11_17_local_g0_1_47128;
  assign net_47129 = seg_11_17_local_g0_2_47129;
  assign net_47131 = seg_11_17_local_g0_4_47131;
  assign net_47132 = seg_11_17_local_g0_5_47132;
  assign net_47135 = seg_11_17_local_g1_0_47135;
  assign net_47136 = seg_11_17_local_g1_1_47136;
  assign net_47137 = seg_11_17_local_g1_2_47137;
  assign net_47138 = seg_11_17_local_g1_3_47138;
  assign net_47141 = seg_11_17_local_g1_6_47141;
  assign net_47143 = seg_11_17_local_g2_0_47143;
  assign net_47145 = seg_11_17_local_g2_2_47145;
  assign net_47156 = seg_11_17_local_g3_5_47156;
  assign net_47250 = seg_11_18_local_g0_0_47250;
  assign net_47251 = seg_11_18_local_g0_1_47251;
  assign net_47252 = seg_11_18_local_g0_2_47252;
  assign net_47255 = seg_11_18_local_g0_5_47255;
  assign net_47256 = seg_11_18_local_g0_6_47256;
  assign net_47257 = seg_11_18_local_g0_7_47257;
  assign net_47260 = seg_11_18_local_g1_2_47260;
  assign net_47263 = seg_11_18_local_g1_5_47263;
  assign net_47264 = seg_11_18_local_g1_6_47264;
  assign net_47265 = seg_11_18_local_g1_7_47265;
  assign net_47266 = seg_11_18_local_g2_0_47266;
  assign net_47268 = seg_11_18_local_g2_2_47268;
  assign net_47277 = seg_11_18_local_g3_3_47277;
  assign net_47278 = seg_11_18_local_g3_4_47278;
  assign net_47280 = seg_11_18_local_g3_6_47280;
  assign net_47382 = seg_11_19_local_g1_1_47382;
  assign net_48952 = seg_12_1_local_g0_2_48952;
  assign net_48954 = seg_12_1_local_g0_4_48954;
  assign net_48959 = seg_12_1_local_g1_1_48959;
  assign net_48967 = seg_12_1_local_g2_1_48967;
  assign net_48968 = seg_12_1_local_g2_2_48968;
  assign net_48975 = seg_12_1_local_g3_1_48975;
  assign net_48977 = seg_12_1_local_g3_3_48977;
  assign net_48979 = seg_12_1_local_g3_5_48979;
  assign net_49115 = seg_12_2_local_g0_2_49115;
  assign net_49119 = seg_12_2_local_g0_6_49119;
  assign net_49123 = seg_12_2_local_g1_2_49123;
  assign net_49124 = seg_12_2_local_g1_3_49124;
  assign net_49131 = seg_12_2_local_g2_2_49131;
  assign net_49134 = seg_12_2_local_g2_5_49134;
  assign net_49236 = seg_12_3_local_g0_0_49236;
  assign net_49238 = seg_12_3_local_g0_2_49238;
  assign net_49239 = seg_12_3_local_g0_3_49239;
  assign net_49240 = seg_12_3_local_g0_4_49240;
  assign net_49241 = seg_12_3_local_g0_5_49241;
  assign net_49246 = seg_12_3_local_g1_2_49246;
  assign net_49256 = seg_12_3_local_g2_4_49256;
  assign net_49257 = seg_12_3_local_g2_5_49257;
  assign net_49258 = seg_12_3_local_g2_6_49258;
  assign net_49266 = seg_12_3_local_g3_6_49266;
  assign net_49363 = seg_12_4_local_g0_4_49363;
  assign net_49365 = seg_12_4_local_g0_6_49365;
  assign net_49366 = seg_12_4_local_g0_7_49366;
  assign net_49367 = seg_12_4_local_g1_0_49367;
  assign net_49371 = seg_12_4_local_g1_4_49371;
  assign net_49373 = seg_12_4_local_g1_6_49373;
  assign net_49375 = seg_12_4_local_g2_0_49375;
  assign net_49378 = seg_12_4_local_g2_3_49378;
  assign net_49379 = seg_12_4_local_g2_4_49379;
  assign net_49380 = seg_12_4_local_g2_5_49380;
  assign net_49383 = seg_12_4_local_g3_0_49383;
  assign net_49384 = seg_12_4_local_g3_1_49384;
  assign net_49385 = seg_12_4_local_g3_2_49385;
  assign net_49386 = seg_12_4_local_g3_3_49386;
  assign net_49388 = seg_12_4_local_g3_5_49388;
  assign net_49390 = seg_12_4_local_g3_7_49390;
  assign net_49493 = seg_12_5_local_g1_3_49493;
  assign net_49494 = seg_12_5_local_g1_4_49494;
  assign net_49495 = seg_12_5_local_g1_5_49495;
  assign net_49511 = seg_12_5_local_g3_5_49511;
  assign net_49608 = seg_12_6_local_g0_3_49608;
  assign net_49610 = seg_12_6_local_g0_5_49610;
  assign net_49616 = seg_12_6_local_g1_3_49616;
  assign net_49617 = seg_12_6_local_g1_4_49617;
  assign net_49620 = seg_12_6_local_g1_7_49620;
  assign net_49623 = seg_12_6_local_g2_2_49623;
  assign net_49629 = seg_12_6_local_g3_0_49629;
  assign net_49630 = seg_12_6_local_g3_1_49630;
  assign net_49636 = seg_12_6_local_g3_7_49636;
  assign net_49737 = seg_12_7_local_g1_1_49737;
  assign net_49739 = seg_12_7_local_g1_3_49739;
  assign net_49741 = seg_12_7_local_g1_5_49741;
  assign net_49742 = seg_12_7_local_g1_6_49742;
  assign net_49744 = seg_12_7_local_g2_0_49744;
  assign net_49745 = seg_12_7_local_g2_1_49745;
  assign net_49750 = seg_12_7_local_g2_6_49750;
  assign net_49752 = seg_12_7_local_g3_0_49752;
  assign net_49755 = seg_12_7_local_g3_3_49755;
  assign net_49855 = seg_12_8_local_g0_4_49855;
  assign net_49857 = seg_12_8_local_g0_6_49857;
  assign net_49859 = seg_12_8_local_g1_0_49859;
  assign net_49861 = seg_12_8_local_g1_2_49861;
  assign net_49985 = seg_12_9_local_g1_3_49985;
  assign net_49993 = seg_12_9_local_g2_3_49993;
  assign net_49998 = seg_12_9_local_g3_0_49998;
  assign net_5 = seg_23_9_glb_netwk_0_5;
  assign net_50001 = seg_12_9_local_g3_3_50001;
  assign net_50097 = seg_12_10_local_g0_0_50097;
  assign net_50100 = seg_12_10_local_g0_3_50100;
  assign net_50101 = seg_12_10_local_g0_4_50101;
  assign net_50108 = seg_12_10_local_g1_3_50108;
  assign net_50110 = seg_12_10_local_g1_5_50110;
  assign net_50122 = seg_12_10_local_g3_1_50122;
  assign net_50222 = seg_12_11_local_g0_2_50222;
  assign net_50224 = seg_12_11_local_g0_4_50224;
  assign net_50227 = seg_12_11_local_g0_7_50227;
  assign net_50231 = seg_12_11_local_g1_3_50231;
  assign net_50233 = seg_12_11_local_g1_5_50233;
  assign net_50235 = seg_12_11_local_g1_7_50235;
  assign net_50345 = seg_12_12_local_g0_2_50345;
  assign net_50353 = seg_12_12_local_g1_2_50353;
  assign net_50355 = seg_12_12_local_g1_4_50355;
  assign net_50362 = seg_12_12_local_g2_3_50362;
  assign net_50363 = seg_12_12_local_g2_4_50363;
  assign net_50368 = seg_12_12_local_g3_1_50368;
  assign net_50372 = seg_12_12_local_g3_5_50372;
  assign net_50466 = seg_12_13_local_g0_0_50466;
  assign net_50472 = seg_12_13_local_g0_6_50472;
  assign net_50475 = seg_12_13_local_g1_1_50475;
  assign net_50476 = seg_12_13_local_g1_2_50476;
  assign net_50477 = seg_12_13_local_g1_3_50477;
  assign net_50492 = seg_12_13_local_g3_2_50492;
  assign net_50494 = seg_12_13_local_g3_4_50494;
  assign net_50590 = seg_12_14_local_g0_1_50590;
  assign net_50598 = seg_12_14_local_g1_1_50598;
  assign net_50599 = seg_12_14_local_g1_2_50599;
  assign net_50600 = seg_12_14_local_g1_3_50600;
  assign net_50602 = seg_12_14_local_g1_5_50602;
  assign net_50606 = seg_12_14_local_g2_1_50606;
  assign net_50609 = seg_12_14_local_g2_4_50609;
  assign net_50612 = seg_12_14_local_g2_7_50612;
  assign net_50614 = seg_12_14_local_g3_1_50614;
  assign net_50616 = seg_12_14_local_g3_3_50616;
  assign net_50617 = seg_12_14_local_g3_4_50617;
  assign net_50619 = seg_12_14_local_g3_6_50619;
  assign net_50714 = seg_12_15_local_g0_2_50714;
  assign net_50715 = seg_12_15_local_g0_3_50715;
  assign net_50723 = seg_12_15_local_g1_3_50723;
  assign net_50724 = seg_12_15_local_g1_4_50724;
  assign net_50731 = seg_12_15_local_g2_3_50731;
  assign net_50734 = seg_12_15_local_g2_6_50734;
  assign net_50739 = seg_12_15_local_g3_3_50739;
  assign net_50740 = seg_12_15_local_g3_4_50740;
  assign net_50742 = seg_12_15_local_g3_6_50742;
  assign net_50835 = seg_12_16_local_g0_0_50835;
  assign net_50836 = seg_12_16_local_g0_1_50836;
  assign net_50837 = seg_12_16_local_g0_2_50837;
  assign net_50838 = seg_12_16_local_g0_3_50838;
  assign net_50839 = seg_12_16_local_g0_4_50839;
  assign net_50840 = seg_12_16_local_g0_5_50840;
  assign net_50841 = seg_12_16_local_g0_6_50841;
  assign net_50842 = seg_12_16_local_g0_7_50842;
  assign net_50844 = seg_12_16_local_g1_1_50844;
  assign net_50846 = seg_12_16_local_g1_3_50846;
  assign net_50847 = seg_12_16_local_g1_4_50847;
  assign net_50848 = seg_12_16_local_g1_5_50848;
  assign net_50849 = seg_12_16_local_g1_6_50849;
  assign net_50850 = seg_12_16_local_g1_7_50850;
  assign net_50856 = seg_12_16_local_g2_5_50856;
  assign net_50857 = seg_12_16_local_g2_6_50857;
  assign net_50858 = seg_12_16_local_g2_7_50858;
  assign net_50864 = seg_12_16_local_g3_5_50864;
  assign net_50866 = seg_12_16_local_g3_7_50866;
  assign net_50959 = seg_12_17_local_g0_1_50959;
  assign net_50966 = seg_12_17_local_g1_0_50966;
  assign net_50971 = seg_12_17_local_g1_5_50971;
  assign net_50978 = seg_12_17_local_g2_4_50978;
  assign net_51082 = seg_12_18_local_g0_1_51082;
  assign net_51092 = seg_12_18_local_g1_3_51092;
  assign net_51093 = seg_12_18_local_g1_4_51093;
  assign net_5117 = seg_0_24_local_g0_2_5117;
  assign net_5118 = seg_0_24_local_g0_3_5118;
  assign net_5120 = seg_0_24_local_g0_5_5120;
  assign net_51218 = seg_12_19_local_g1_6_51218;
  assign net_5122 = seg_0_24_local_g0_7_5122;
  assign net_5123 = seg_0_24_local_g1_0_5123;
  assign net_51231 = seg_12_19_local_g3_3_51231;
  assign net_5125 = seg_0_24_local_g1_2_5125;
  assign net_5126 = seg_0_24_local_g1_3_5126;
  assign net_5127 = seg_0_24_local_g1_4_5127;
  assign net_5128 = seg_0_24_local_g1_5_5128;
  assign net_5133 = seg_0_24_local_g2_2_5133;
  assign net_5134 = seg_0_24_local_g2_3_5134;
  assign net_5140 = seg_0_24_local_g3_1_5140;
  assign net_5141 = seg_0_24_local_g3_2_5141;
  assign net_5142 = seg_0_24_local_g3_3_5142;
  assign net_5144 = seg_0_24_local_g3_5_5144;
  assign net_5146 = seg_0_24_local_g3_7_5146;
  assign net_52784 = seg_13_1_local_g0_3_52784;
  assign net_52785 = seg_13_1_local_g0_4_52785;
  assign net_52791 = seg_13_1_local_g1_2_52791;
  assign net_52792 = seg_13_1_local_g1_3_52792;
  assign net_52793 = seg_13_1_local_g1_4_52793;
  assign net_52948 = seg_13_2_local_g0_4_52948;
  assign net_52952 = seg_13_2_local_g1_0_52952;
  assign net_52954 = seg_13_2_local_g1_2_52954;
  assign net_52955 = seg_13_2_local_g1_3_52955;
  assign net_52959 = seg_13_2_local_g1_7_52959;
  assign net_52963 = seg_13_2_local_g2_3_52963;
  assign net_52970 = seg_13_2_local_g3_2_52970;
  assign net_52971 = seg_13_2_local_g3_3_52971;
  assign net_53067 = seg_13_3_local_g0_0_53067;
  assign net_53068 = seg_13_3_local_g0_1_53068;
  assign net_53070 = seg_13_3_local_g0_3_53070;
  assign net_53073 = seg_13_3_local_g0_6_53073;
  assign net_53074 = seg_13_3_local_g0_7_53074;
  assign net_53080 = seg_13_3_local_g1_5_53080;
  assign net_53083 = seg_13_3_local_g2_0_53083;
  assign net_53087 = seg_13_3_local_g2_4_53087;
  assign net_53088 = seg_13_3_local_g2_5_53088;
  assign net_53092 = seg_13_3_local_g3_1_53092;
  assign net_53093 = seg_13_3_local_g3_2_53093;
  assign net_53192 = seg_13_4_local_g0_2_53192;
  assign net_53193 = seg_13_4_local_g0_3_53193;
  assign net_53194 = seg_13_4_local_g0_4_53194;
  assign net_53195 = seg_13_4_local_g0_5_53195;
  assign net_53198 = seg_13_4_local_g1_0_53198;
  assign net_53199 = seg_13_4_local_g1_1_53199;
  assign net_53200 = seg_13_4_local_g1_2_53200;
  assign net_53201 = seg_13_4_local_g1_3_53201;
  assign net_53203 = seg_13_4_local_g1_5_53203;
  assign net_53206 = seg_13_4_local_g2_0_53206;
  assign net_53207 = seg_13_4_local_g2_1_53207;
  assign net_53210 = seg_13_4_local_g2_4_53210;
  assign net_53211 = seg_13_4_local_g2_5_53211;
  assign net_53217 = seg_13_4_local_g3_3_53217;
  assign net_5323 = seg_0_25_local_g0_2_5323;
  assign net_5325 = seg_0_25_local_g0_4_5325;
  assign net_5326 = seg_0_25_local_g0_5_5326;
  assign net_5327 = seg_0_25_local_g0_6_5327;
  assign net_5328 = seg_0_25_local_g0_7_5328;
  assign net_5329 = seg_0_25_local_g1_0_5329;
  assign net_5330 = seg_0_25_local_g1_1_5330;
  assign net_5331 = seg_0_25_local_g1_2_5331;
  assign net_53315 = seg_13_5_local_g0_2_53315;
  assign net_5332 = seg_0_25_local_g1_3_5332;
  assign net_53322 = seg_13_5_local_g1_1_53322;
  assign net_53324 = seg_13_5_local_g1_3_53324;
  assign net_53331 = seg_13_5_local_g2_2_53331;
  assign net_53332 = seg_13_5_local_g2_3_53332;
  assign net_5336 = seg_0_25_local_g1_7_5336;
  assign net_5340 = seg_0_25_local_g2_3_5340;
  assign net_5341 = seg_0_25_local_g2_4_5341;
  assign net_5342 = seg_0_25_local_g2_5_5342;
  assign net_53439 = seg_13_6_local_g0_3_53439;
  assign net_5344 = seg_0_25_local_g2_7_5344;
  assign net_53441 = seg_13_6_local_g0_5_53441;
  assign net_53445 = seg_13_6_local_g1_1_53445;
  assign net_5345 = seg_0_25_local_g3_0_5345;
  assign net_53450 = seg_13_6_local_g1_6_53450;
  assign net_53451 = seg_13_6_local_g1_7_53451;
  assign net_53453 = seg_13_6_local_g2_1_53453;
  assign net_53454 = seg_13_6_local_g2_2_53454;
  assign net_53455 = seg_13_6_local_g2_3_53455;
  assign net_53458 = seg_13_6_local_g2_6_53458;
  assign net_5346 = seg_0_25_local_g3_1_5346;
  assign net_53462 = seg_13_6_local_g3_2_53462;
  assign net_53467 = seg_13_6_local_g3_7_53467;
  assign net_53559 = seg_13_7_local_g0_0_53559;
  assign net_53564 = seg_13_7_local_g0_5_53564;
  assign net_53566 = seg_13_7_local_g0_7_53566;
  assign net_53567 = seg_13_7_local_g1_0_53567;
  assign net_53569 = seg_13_7_local_g1_2_53569;
  assign net_53570 = seg_13_7_local_g1_3_53570;
  assign net_53578 = seg_13_7_local_g2_3_53578;
  assign net_53579 = seg_13_7_local_g2_4_53579;
  assign net_53580 = seg_13_7_local_g2_5_53580;
  assign net_53584 = seg_13_7_local_g3_1_53584;
  assign net_53586 = seg_13_7_local_g3_3_53586;
  assign net_53587 = seg_13_7_local_g3_4_53587;
  assign net_53588 = seg_13_7_local_g3_5_53588;
  assign net_53589 = seg_13_7_local_g3_6_53589;
  assign net_53590 = seg_13_7_local_g3_7_53590;
  assign net_53682 = seg_13_8_local_g0_0_53682;
  assign net_53684 = seg_13_8_local_g0_2_53684;
  assign net_53685 = seg_13_8_local_g0_3_53685;
  assign net_53686 = seg_13_8_local_g0_4_53686;
  assign net_53687 = seg_13_8_local_g0_5_53687;
  assign net_53688 = seg_13_8_local_g0_6_53688;
  assign net_53691 = seg_13_8_local_g1_1_53691;
  assign net_53692 = seg_13_8_local_g1_2_53692;
  assign net_53693 = seg_13_8_local_g1_3_53693;
  assign net_53695 = seg_13_8_local_g1_5_53695;
  assign net_53696 = seg_13_8_local_g1_6_53696;
  assign net_53699 = seg_13_8_local_g2_1_53699;
  assign net_53701 = seg_13_8_local_g2_3_53701;
  assign net_53702 = seg_13_8_local_g2_4_53702;
  assign net_53703 = seg_13_8_local_g2_5_53703;
  assign net_53711 = seg_13_8_local_g3_5_53711;
  assign net_53712 = seg_13_8_local_g3_6_53712;
  assign net_53811 = seg_13_9_local_g0_6_53811;
  assign net_53816 = seg_13_9_local_g1_3_53816;
  assign net_53832 = seg_13_9_local_g3_3_53832;
  assign net_53929 = seg_13_10_local_g0_1_53929;
  assign net_53940 = seg_13_10_local_g1_4_53940;
  assign net_53941 = seg_13_10_local_g1_5_53941;
  assign net_53942 = seg_13_10_local_g1_6_53942;
  assign net_53944 = seg_13_10_local_g2_0_53944;
  assign net_53945 = seg_13_10_local_g2_1_53945;
  assign net_53946 = seg_13_10_local_g2_2_53946;
  assign net_53949 = seg_13_10_local_g2_5_53949;
  assign net_53952 = seg_13_10_local_g3_0_53952;
  assign net_53953 = seg_13_10_local_g3_1_53953;
  assign net_53955 = seg_13_10_local_g3_3_53955;
  assign net_54055 = seg_13_11_local_g0_4_54055;
  assign net_54056 = seg_13_11_local_g0_5_54056;
  assign net_54058 = seg_13_11_local_g0_7_54058;
  assign net_54066 = seg_13_11_local_g1_7_54066;
  assign net_54070 = seg_13_11_local_g2_3_54070;
  assign net_54072 = seg_13_11_local_g2_5_54072;
  assign net_54073 = seg_13_11_local_g2_6_54073;
  assign net_54078 = seg_13_11_local_g3_3_54078;
  assign net_54082 = seg_13_11_local_g3_7_54082;
  assign net_54176 = seg_13_12_local_g0_2_54176;
  assign net_54179 = seg_13_12_local_g0_5_54179;
  assign net_54180 = seg_13_12_local_g0_6_54180;
  assign net_54183 = seg_13_12_local_g1_1_54183;
  assign net_54184 = seg_13_12_local_g1_2_54184;
  assign net_54195 = seg_13_12_local_g2_5_54195;
  assign net_54196 = seg_13_12_local_g2_6_54196;
  assign net_54199 = seg_13_12_local_g3_1_54199;
  assign net_54205 = seg_13_12_local_g3_7_54205;
  assign net_54299 = seg_13_13_local_g0_2_54299;
  assign net_54303 = seg_13_13_local_g0_6_54303;
  assign net_54304 = seg_13_13_local_g0_7_54304;
  assign net_54305 = seg_13_13_local_g1_0_54305;
  assign net_54307 = seg_13_13_local_g1_2_54307;
  assign net_54308 = seg_13_13_local_g1_3_54308;
  assign net_54309 = seg_13_13_local_g1_4_54309;
  assign net_54311 = seg_13_13_local_g1_6_54311;
  assign net_54313 = seg_13_13_local_g2_0_54313;
  assign net_54316 = seg_13_13_local_g2_3_54316;
  assign net_54317 = seg_13_13_local_g2_4_54317;
  assign net_54323 = seg_13_13_local_g3_2_54323;
  assign net_54324 = seg_13_13_local_g3_3_54324;
  assign net_54325 = seg_13_13_local_g3_4_54325;
  assign net_54326 = seg_13_13_local_g3_5_54326;
  assign net_54425 = seg_13_14_local_g0_5_54425;
  assign net_54427 = seg_13_14_local_g0_7_54427;
  assign net_54428 = seg_13_14_local_g1_0_54428;
  assign net_54429 = seg_13_14_local_g1_1_54429;
  assign net_54431 = seg_13_14_local_g1_3_54431;
  assign net_54433 = seg_13_14_local_g1_5_54433;
  assign net_54435 = seg_13_14_local_g1_7_54435;
  assign net_54436 = seg_13_14_local_g2_0_54436;
  assign net_54437 = seg_13_14_local_g2_1_54437;
  assign net_54438 = seg_13_14_local_g2_2_54438;
  assign net_54444 = seg_13_14_local_g3_0_54444;
  assign net_54446 = seg_13_14_local_g3_2_54446;
  assign net_54447 = seg_13_14_local_g3_3_54447;
  assign net_54450 = seg_13_14_local_g3_6_54450;
  assign net_54543 = seg_13_15_local_g0_0_54543;
  assign net_54544 = seg_13_15_local_g0_1_54544;
  assign net_54546 = seg_13_15_local_g0_3_54546;
  assign net_54549 = seg_13_15_local_g0_6_54549;
  assign net_54551 = seg_13_15_local_g1_0_54551;
  assign net_54552 = seg_13_15_local_g1_1_54552;
  assign net_54553 = seg_13_15_local_g1_2_54553;
  assign net_54554 = seg_13_15_local_g1_3_54554;
  assign net_54555 = seg_13_15_local_g1_4_54555;
  assign net_54556 = seg_13_15_local_g1_5_54556;
  assign net_54561 = seg_13_15_local_g2_2_54561;
  assign net_54567 = seg_13_15_local_g3_0_54567;
  assign net_54574 = seg_13_15_local_g3_7_54574;
  assign net_54667 = seg_13_16_local_g0_1_54667;
  assign net_54668 = seg_13_16_local_g0_2_54668;
  assign net_54669 = seg_13_16_local_g0_3_54669;
  assign net_54670 = seg_13_16_local_g0_4_54670;
  assign net_54672 = seg_13_16_local_g0_6_54672;
  assign net_54673 = seg_13_16_local_g0_7_54673;
  assign net_54676 = seg_13_16_local_g1_2_54676;
  assign net_54677 = seg_13_16_local_g1_3_54677;
  assign net_54678 = seg_13_16_local_g1_4_54678;
  assign net_54679 = seg_13_16_local_g1_5_54679;
  assign net_54682 = seg_13_16_local_g2_0_54682;
  assign net_54685 = seg_13_16_local_g2_3_54685;
  assign net_54694 = seg_13_16_local_g3_4_54694;
  assign net_54695 = seg_13_16_local_g3_5_54695;
  assign net_54696 = seg_13_16_local_g3_6_54696;
  assign net_54789 = seg_13_17_local_g0_0_54789;
  assign net_54790 = seg_13_17_local_g0_1_54790;
  assign net_54793 = seg_13_17_local_g0_4_54793;
  assign net_54796 = seg_13_17_local_g0_7_54796;
  assign net_54800 = seg_13_17_local_g1_3_54800;
  assign net_54803 = seg_13_17_local_g1_6_54803;
  assign net_54804 = seg_13_17_local_g1_7_54804;
  assign net_54816 = seg_13_17_local_g3_3_54816;
  assign net_54912 = seg_13_18_local_g0_0_54912;
  assign net_54913 = seg_13_18_local_g0_1_54913;
  assign net_54915 = seg_13_18_local_g0_3_54915;
  assign net_54916 = seg_13_18_local_g0_4_54916;
  assign net_54917 = seg_13_18_local_g0_5_54917;
  assign net_54919 = seg_13_18_local_g0_7_54919;
  assign net_54920 = seg_13_18_local_g1_0_54920;
  assign net_54923 = seg_13_18_local_g1_3_54923;
  assign net_54924 = seg_13_18_local_g1_4_54924;
  assign net_54925 = seg_13_18_local_g1_5_54925;
  assign net_54926 = seg_13_18_local_g1_6_54926;
  assign net_54927 = seg_13_18_local_g1_7_54927;
  assign net_54928 = seg_13_18_local_g2_0_54928;
  assign net_54929 = seg_13_18_local_g2_1_54929;
  assign net_54930 = seg_13_18_local_g2_2_54930;
  assign net_54931 = seg_13_18_local_g2_3_54931;
  assign net_54933 = seg_13_18_local_g2_5_54933;
  assign net_54935 = seg_13_18_local_g2_7_54935;
  assign net_54936 = seg_13_18_local_g3_0_54936;
  assign net_54938 = seg_13_18_local_g3_2_54938;
  assign net_54939 = seg_13_18_local_g3_3_54939;
  assign net_54941 = seg_13_18_local_g3_5_54941;
  assign net_54942 = seg_13_18_local_g3_6_54942;
  assign net_55036 = seg_13_19_local_g0_1_55036;
  assign net_55039 = seg_13_19_local_g0_4_55039;
  assign net_55044 = seg_13_19_local_g1_1_55044;
  assign net_55046 = seg_13_19_local_g1_3_55046;
  assign net_55049 = seg_13_19_local_g1_6_55049;
  assign net_56527 = seg_13_31_local_g0_3_56527;
  assign net_56533 = seg_13_31_local_g1_1_56533;
  assign net_56614 = seg_14_1_local_g0_3_56614;
  assign net_56627 = seg_14_1_local_g2_0_56627;
  assign net_56774 = seg_14_2_local_g0_0_56774;
  assign net_56776 = seg_14_2_local_g0_2_56776;
  assign net_56779 = seg_14_2_local_g0_5_56779;
  assign net_56783 = seg_14_2_local_g1_1_56783;
  assign net_56785 = seg_14_2_local_g1_3_56785;
  assign net_56788 = seg_14_2_local_g1_6_56788;
  assign net_56900 = seg_14_3_local_g0_3_56900;
  assign net_56907 = seg_14_3_local_g1_2_56907;
  assign net_57020 = seg_14_4_local_g0_0_57020;
  assign net_57026 = seg_14_4_local_g0_6_57026;
  assign net_57032 = seg_14_4_local_g1_4_57032;
  assign net_57035 = seg_14_4_local_g1_7_57035;
  assign net_57040 = seg_14_4_local_g2_4_57040;
  assign net_57043 = seg_14_4_local_g2_7_57043;
  assign net_57045 = seg_14_4_local_g3_1_57045;
  assign net_57048 = seg_14_4_local_g3_4_57048;
  assign net_57051 = seg_14_4_local_g3_7_57051;
  assign net_57143 = seg_14_5_local_g0_0_57143;
  assign net_57145 = seg_14_5_local_g0_2_57145;
  assign net_57146 = seg_14_5_local_g0_3_57146;
  assign net_57152 = seg_14_5_local_g1_1_57152;
  assign net_57155 = seg_14_5_local_g1_4_57155;
  assign net_57156 = seg_14_5_local_g1_5_57156;
  assign net_57159 = seg_14_5_local_g2_0_57159;
  assign net_57160 = seg_14_5_local_g2_1_57160;
  assign net_57162 = seg_14_5_local_g2_3_57162;
  assign net_57163 = seg_14_5_local_g2_4_57163;
  assign net_57165 = seg_14_5_local_g2_6_57165;
  assign net_57166 = seg_14_5_local_g2_7_57166;
  assign net_57168 = seg_14_5_local_g3_1_57168;
  assign net_57170 = seg_14_5_local_g3_3_57170;
  assign net_57172 = seg_14_5_local_g3_5_57172;
  assign net_57173 = seg_14_5_local_g3_6_57173;
  assign net_57174 = seg_14_5_local_g3_7_57174;
  assign net_57266 = seg_14_6_local_g0_0_57266;
  assign net_57269 = seg_14_6_local_g0_3_57269;
  assign net_57270 = seg_14_6_local_g0_4_57270;
  assign net_57273 = seg_14_6_local_g0_7_57273;
  assign net_57275 = seg_14_6_local_g1_1_57275;
  assign net_57276 = seg_14_6_local_g1_2_57276;
  assign net_57277 = seg_14_6_local_g1_3_57277;
  assign net_57278 = seg_14_6_local_g1_4_57278;
  assign net_57279 = seg_14_6_local_g1_5_57279;
  assign net_57282 = seg_14_6_local_g2_0_57282;
  assign net_57288 = seg_14_6_local_g2_6_57288;
  assign net_57290 = seg_14_6_local_g3_0_57290;
  assign net_57294 = seg_14_6_local_g3_4_57294;
  assign net_57295 = seg_14_6_local_g3_5_57295;
  assign net_57296 = seg_14_6_local_g3_6_57296;
  assign net_57396 = seg_14_7_local_g0_7_57396;
  assign net_57402 = seg_14_7_local_g1_5_57402;
  assign net_57404 = seg_14_7_local_g1_7_57404;
  assign net_57407 = seg_14_7_local_g2_2_57407;
  assign net_57416 = seg_14_7_local_g3_3_57416;
  assign net_57512 = seg_14_8_local_g0_0_57512;
  assign net_57513 = seg_14_8_local_g0_1_57513;
  assign net_57517 = seg_14_8_local_g0_5_57517;
  assign net_57521 = seg_14_8_local_g1_1_57521;
  assign net_57523 = seg_14_8_local_g1_3_57523;
  assign net_57524 = seg_14_8_local_g1_4_57524;
  assign net_57525 = seg_14_8_local_g1_5_57525;
  assign net_57528 = seg_14_8_local_g2_0_57528;
  assign net_57536 = seg_14_8_local_g3_0_57536;
  assign net_57538 = seg_14_8_local_g3_2_57538;
  assign net_57541 = seg_14_8_local_g3_5_57541;
  assign net_57635 = seg_14_9_local_g0_0_57635;
  assign net_57636 = seg_14_9_local_g0_1_57636;
  assign net_57637 = seg_14_9_local_g0_2_57637;
  assign net_57639 = seg_14_9_local_g0_4_57639;
  assign net_57643 = seg_14_9_local_g1_0_57643;
  assign net_57644 = seg_14_9_local_g1_1_57644;
  assign net_57646 = seg_14_9_local_g1_3_57646;
  assign net_57759 = seg_14_10_local_g0_1_57759;
  assign net_57760 = seg_14_10_local_g0_2_57760;
  assign net_57771 = seg_14_10_local_g1_5_57771;
  assign net_57773 = seg_14_10_local_g1_7_57773;
  assign net_57774 = seg_14_10_local_g2_0_57774;
  assign net_57778 = seg_14_10_local_g2_4_57778;
  assign net_57781 = seg_14_10_local_g2_7_57781;
  assign net_57782 = seg_14_10_local_g3_0_57782;
  assign net_57786 = seg_14_10_local_g3_4_57786;
  assign net_57883 = seg_14_11_local_g0_2_57883;
  assign net_57884 = seg_14_11_local_g0_3_57884;
  assign net_57890 = seg_14_11_local_g1_1_57890;
  assign net_57893 = seg_14_11_local_g1_4_57893;
  assign net_57896 = seg_14_11_local_g1_7_57896;
  assign net_58012 = seg_14_12_local_g1_0_58012;
  assign net_58131 = seg_14_13_local_g0_4_58131;
  assign net_58133 = seg_14_13_local_g0_6_58133;
  assign net_58139 = seg_14_13_local_g1_4_58139;
  assign net_58143 = seg_14_13_local_g2_0_58143;
  assign net_58144 = seg_14_13_local_g2_1_58144;
  assign net_58145 = seg_14_13_local_g2_2_58145;
  assign net_58147 = seg_14_13_local_g2_4_58147;
  assign net_58151 = seg_14_13_local_g3_0_58151;
  assign net_58152 = seg_14_13_local_g3_1_58152;
  assign net_58154 = seg_14_13_local_g3_3_58154;
  assign net_58155 = seg_14_13_local_g3_4_58155;
  assign net_58250 = seg_14_14_local_g0_0_58250;
  assign net_58251 = seg_14_14_local_g0_1_58251;
  assign net_58253 = seg_14_14_local_g0_3_58253;
  assign net_58254 = seg_14_14_local_g0_4_58254;
  assign net_58264 = seg_14_14_local_g1_6_58264;
  assign net_58268 = seg_14_14_local_g2_2_58268;
  assign net_58270 = seg_14_14_local_g2_4_58270;
  assign net_58273 = seg_14_14_local_g2_7_58273;
  assign net_58274 = seg_14_14_local_g3_0_58274;
  assign net_58275 = seg_14_14_local_g3_1_58275;
  assign net_58373 = seg_14_15_local_g0_0_58373;
  assign net_58375 = seg_14_15_local_g0_2_58375;
  assign net_58378 = seg_14_15_local_g0_5_58378;
  assign net_58380 = seg_14_15_local_g0_7_58380;
  assign net_58385 = seg_14_15_local_g1_4_58385;
  assign net_58386 = seg_14_15_local_g1_5_58386;
  assign net_58387 = seg_14_15_local_g1_6_58387;
  assign net_58388 = seg_14_15_local_g1_7_58388;
  assign net_58393 = seg_14_15_local_g2_4_58393;
  assign net_58396 = seg_14_15_local_g2_7_58396;
  assign net_58496 = seg_14_16_local_g0_0_58496;
  assign net_58499 = seg_14_16_local_g0_3_58499;
  assign net_58500 = seg_14_16_local_g0_4_58500;
  assign net_58501 = seg_14_16_local_g0_5_58501;
  assign net_58503 = seg_14_16_local_g0_7_58503;
  assign net_58504 = seg_14_16_local_g1_0_58504;
  assign net_58506 = seg_14_16_local_g1_2_58506;
  assign net_58507 = seg_14_16_local_g1_3_58507;
  assign net_58509 = seg_14_16_local_g1_5_58509;
  assign net_58510 = seg_14_16_local_g1_6_58510;
  assign net_58511 = seg_14_16_local_g1_7_58511;
  assign net_58514 = seg_14_16_local_g2_2_58514;
  assign net_58516 = seg_14_16_local_g2_4_58516;
  assign net_58522 = seg_14_16_local_g3_2_58522;
  assign net_58527 = seg_14_16_local_g3_7_58527;
  assign net_58620 = seg_14_17_local_g0_1_58620;
  assign net_58621 = seg_14_17_local_g0_2_58621;
  assign net_58626 = seg_14_17_local_g0_7_58626;
  assign net_58630 = seg_14_17_local_g1_3_58630;
  assign net_58633 = seg_14_17_local_g1_6_58633;
  assign net_58646 = seg_14_17_local_g3_3_58646;
  assign net_58742 = seg_14_18_local_g0_0_58742;
  assign net_58743 = seg_14_18_local_g0_1_58743;
  assign net_58745 = seg_14_18_local_g0_3_58745;
  assign net_58747 = seg_14_18_local_g0_5_58747;
  assign net_58748 = seg_14_18_local_g0_6_58748;
  assign net_58750 = seg_14_18_local_g1_0_58750;
  assign net_58751 = seg_14_18_local_g1_1_58751;
  assign net_58752 = seg_14_18_local_g1_2_58752;
  assign net_58753 = seg_14_18_local_g1_3_58753;
  assign net_58754 = seg_14_18_local_g1_4_58754;
  assign net_58756 = seg_14_18_local_g1_6_58756;
  assign net_58761 = seg_14_18_local_g2_3_58761;
  assign net_58764 = seg_14_18_local_g2_6_58764;
  assign net_58765 = seg_14_18_local_g2_7_58765;
  assign net_58768 = seg_14_18_local_g3_2_58768;
  assign net_58769 = seg_14_18_local_g3_3_58769;
  assign net_58770 = seg_14_18_local_g3_4_58770;
  assign net_58883 = seg_14_19_local_g2_2_58883;
  assign net_58884 = seg_14_19_local_g2_3_58884;
  assign net_58889 = seg_14_19_local_g3_0_58889;
  assign net_58892 = seg_14_19_local_g3_3_58892;
  assign net_58896 = seg_14_19_local_g3_7_58896;
  assign net_6 = seg_20_12_glb_netwk_1_6;
  assign net_60627 = seg_15_2_local_g2_7_60627;
  assign net_60729 = seg_15_3_local_g0_2_60729;
  assign net_60731 = seg_15_3_local_g0_4_60731;
  assign net_60850 = seg_15_4_local_g0_0_60850;
  assign net_60852 = seg_15_4_local_g0_2_60852;
  assign net_60860 = seg_15_4_local_g1_2_60860;
  assign net_60866 = seg_15_4_local_g2_0_60866;
  assign net_60870 = seg_15_4_local_g2_4_60870;
  assign net_60874 = seg_15_4_local_g3_0_60874;
  assign net_60876 = seg_15_4_local_g3_2_60876;
  assign net_60878 = seg_15_4_local_g3_4_60878;
  assign net_60880 = seg_15_4_local_g3_6_60880;
  assign net_60973 = seg_15_5_local_g0_0_60973;
  assign net_60978 = seg_15_5_local_g0_5_60978;
  assign net_60982 = seg_15_5_local_g1_1_60982;
  assign net_60983 = seg_15_5_local_g1_2_60983;
  assign net_60988 = seg_15_5_local_g1_7_60988;
  assign net_60991 = seg_15_5_local_g2_2_60991;
  assign net_60993 = seg_15_5_local_g2_4_60993;
  assign net_60998 = seg_15_5_local_g3_1_60998;
  assign net_61001 = seg_15_5_local_g3_4_61001;
  assign net_61096 = seg_15_6_local_g0_0_61096;
  assign net_61097 = seg_15_6_local_g0_1_61097;
  assign net_61098 = seg_15_6_local_g0_2_61098;
  assign net_61099 = seg_15_6_local_g0_3_61099;
  assign net_61100 = seg_15_6_local_g0_4_61100;
  assign net_61102 = seg_15_6_local_g0_6_61102;
  assign net_61104 = seg_15_6_local_g1_0_61104;
  assign net_61106 = seg_15_6_local_g1_2_61106;
  assign net_61107 = seg_15_6_local_g1_3_61107;
  assign net_61108 = seg_15_6_local_g1_4_61108;
  assign net_61109 = seg_15_6_local_g1_5_61109;
  assign net_61111 = seg_15_6_local_g1_7_61111;
  assign net_61112 = seg_15_6_local_g2_0_61112;
  assign net_61114 = seg_15_6_local_g2_2_61114;
  assign net_61115 = seg_15_6_local_g2_3_61115;
  assign net_61116 = seg_15_6_local_g2_4_61116;
  assign net_61117 = seg_15_6_local_g2_5_61117;
  assign net_61118 = seg_15_6_local_g2_6_61118;
  assign net_61121 = seg_15_6_local_g3_1_61121;
  assign net_61122 = seg_15_6_local_g3_2_61122;
  assign net_61123 = seg_15_6_local_g3_3_61123;
  assign net_61124 = seg_15_6_local_g3_4_61124;
  assign net_61125 = seg_15_6_local_g3_5_61125;
  assign net_61127 = seg_15_6_local_g3_7_61127;
  assign net_61234 = seg_15_7_local_g1_7_61234;
  assign net_61241 = seg_15_7_local_g2_6_61241;
  assign net_61242 = seg_15_7_local_g2_7_61242;
  assign net_61246 = seg_15_7_local_g3_3_61246;
  assign net_61345 = seg_15_8_local_g0_3_61345;
  assign net_61347 = seg_15_8_local_g0_5_61347;
  assign net_61355 = seg_15_8_local_g1_5_61355;
  assign net_61366 = seg_15_8_local_g3_0_61366;
  assign net_61468 = seg_15_9_local_g0_3_61468;
  assign net_61469 = seg_15_9_local_g0_4_61469;
  assign net_61475 = seg_15_9_local_g1_2_61475;
  assign net_61476 = seg_15_9_local_g1_3_61476;
  assign net_61485 = seg_15_9_local_g2_4_61485;
  assign net_61492 = seg_15_9_local_g3_3_61492;
  assign net_61496 = seg_15_9_local_g3_7_61496;
  assign net_61588 = seg_15_10_local_g0_0_61588;
  assign net_61594 = seg_15_10_local_g0_6_61594;
  assign net_61596 = seg_15_10_local_g1_0_61596;
  assign net_61597 = seg_15_10_local_g1_1_61597;
  assign net_61602 = seg_15_10_local_g1_6_61602;
  assign net_61606 = seg_15_10_local_g2_2_61606;
  assign net_61607 = seg_15_10_local_g2_3_61607;
  assign net_61610 = seg_15_10_local_g2_6_61610;
  assign net_61614 = seg_15_10_local_g3_2_61614;
  assign net_61713 = seg_15_11_local_g0_2_61713;
  assign net_61714 = seg_15_11_local_g0_3_61714;
  assign net_61720 = seg_15_11_local_g1_1_61720;
  assign net_61723 = seg_15_11_local_g1_4_61723;
  assign net_61724 = seg_15_11_local_g1_5_61724;
  assign net_61725 = seg_15_11_local_g1_6_61725;
  assign net_61731 = seg_15_11_local_g2_4_61731;
  assign net_61733 = seg_15_11_local_g2_6_61733;
  assign net_61734 = seg_15_11_local_g2_7_61734;
  assign net_61736 = seg_15_11_local_g3_1_61736;
  assign net_61737 = seg_15_11_local_g3_2_61737;
  assign net_61742 = seg_15_11_local_g3_7_61742;
  assign net_61841 = seg_15_12_local_g0_7_61841;
  assign net_61843 = seg_15_12_local_g1_1_61843;
  assign net_61849 = seg_15_12_local_g1_7_61849;
  assign net_61851 = seg_15_12_local_g2_1_61851;
  assign net_61852 = seg_15_12_local_g2_2_61852;
  assign net_61854 = seg_15_12_local_g2_4_61854;
  assign net_61857 = seg_15_12_local_g2_7_61857;
  assign net_61864 = seg_15_12_local_g3_6_61864;
  assign net_61865 = seg_15_12_local_g3_7_61865;
  assign net_61962 = seg_15_13_local_g0_5_61962;
  assign net_61968 = seg_15_13_local_g1_3_61968;
  assign net_61975 = seg_15_13_local_g2_2_61975;
  assign net_61976 = seg_15_13_local_g2_3_61976;
  assign net_61982 = seg_15_13_local_g3_1_61982;
  assign net_61985 = seg_15_13_local_g3_4_61985;
  assign net_61986 = seg_15_13_local_g3_5_61986;
  assign net_61987 = seg_15_13_local_g3_6_61987;
  assign net_62081 = seg_15_14_local_g0_1_62081;
  assign net_62082 = seg_15_14_local_g0_2_62082;
  assign net_62083 = seg_15_14_local_g0_3_62083;
  assign net_62085 = seg_15_14_local_g0_5_62085;
  assign net_62090 = seg_15_14_local_g1_2_62090;
  assign net_62091 = seg_15_14_local_g1_3_62091;
  assign net_62092 = seg_15_14_local_g1_4_62092;
  assign net_62093 = seg_15_14_local_g1_5_62093;
  assign net_62096 = seg_15_14_local_g2_0_62096;
  assign net_62097 = seg_15_14_local_g2_1_62097;
  assign net_62107 = seg_15_14_local_g3_3_62107;
  assign net_62109 = seg_15_14_local_g3_5_62109;
  assign net_62212 = seg_15_15_local_g1_1_62212;
  assign net_62213 = seg_15_15_local_g1_2_62213;
  assign net_62214 = seg_15_15_local_g1_3_62214;
  assign net_62228 = seg_15_15_local_g3_1_62228;
  assign net_62232 = seg_15_15_local_g3_5_62232;
  assign net_62233 = seg_15_15_local_g3_6_62233;
  assign net_62326 = seg_15_16_local_g0_0_62326;
  assign net_62327 = seg_15_16_local_g0_1_62327;
  assign net_62331 = seg_15_16_local_g0_5_62331;
  assign net_62333 = seg_15_16_local_g0_7_62333;
  assign net_62335 = seg_15_16_local_g1_1_62335;
  assign net_62337 = seg_15_16_local_g1_3_62337;
  assign net_62342 = seg_15_16_local_g2_0_62342;
  assign net_62345 = seg_15_16_local_g2_3_62345;
  assign net_62347 = seg_15_16_local_g2_5_62347;
  assign net_62348 = seg_15_16_local_g2_6_62348;
  assign net_62351 = seg_15_16_local_g3_1_62351;
  assign net_62352 = seg_15_16_local_g3_2_62352;
  assign net_62353 = seg_15_16_local_g3_3_62353;
  assign net_62355 = seg_15_16_local_g3_5_62355;
  assign net_62356 = seg_15_16_local_g3_6_62356;
  assign net_62449 = seg_15_17_local_g0_0_62449;
  assign net_62466 = seg_15_17_local_g2_1_62466;
  assign net_62467 = seg_15_17_local_g2_2_62467;
  assign net_62468 = seg_15_17_local_g2_3_62468;
  assign net_62470 = seg_15_17_local_g2_5_62470;
  assign net_62480 = seg_15_17_local_g3_7_62480;
  assign net_62575 = seg_15_18_local_g0_3_62575;
  assign net_62582 = seg_15_18_local_g1_2_62582;
  assign net_62583 = seg_15_18_local_g1_3_62583;
  assign net_62592 = seg_15_18_local_g2_4_62592;
  assign net_62597 = seg_15_18_local_g3_1_62597;
  assign net_64225 = seg_16_0_local_g1_3_64225;
  assign net_64440 = seg_16_2_local_g0_5_64440;
  assign net_64560 = seg_16_3_local_g0_2_64560;
  assign net_64564 = seg_16_3_local_g0_6_64564;
  assign net_64568 = seg_16_3_local_g1_2_64568;
  assign net_64569 = seg_16_3_local_g1_3_64569;
  assign net_64580 = seg_16_3_local_g2_6_64580;
  assign net_64585 = seg_16_3_local_g3_3_64585;
  assign net_64586 = seg_16_3_local_g3_4_64586;
  assign net_64685 = seg_16_4_local_g0_4_64685;
  assign net_64688 = seg_16_4_local_g0_7_64688;
  assign net_64692 = seg_16_4_local_g1_3_64692;
  assign net_64693 = seg_16_4_local_g1_4_64693;
  assign net_64695 = seg_16_4_local_g1_6_64695;
  assign net_64696 = seg_16_4_local_g1_7_64696;
  assign net_64697 = seg_16_4_local_g2_0_64697;
  assign net_64698 = seg_16_4_local_g2_1_64698;
  assign net_64699 = seg_16_4_local_g2_2_64699;
  assign net_64700 = seg_16_4_local_g2_3_64700;
  assign net_64701 = seg_16_4_local_g2_4_64701;
  assign net_64702 = seg_16_4_local_g2_5_64702;
  assign net_64703 = seg_16_4_local_g2_6_64703;
  assign net_64705 = seg_16_4_local_g3_0_64705;
  assign net_64711 = seg_16_4_local_g3_6_64711;
  assign net_64712 = seg_16_4_local_g3_7_64712;
  assign net_64805 = seg_16_5_local_g0_1_64805;
  assign net_64812 = seg_16_5_local_g1_0_64812;
  assign net_64817 = seg_16_5_local_g1_5_64817;
  assign net_64820 = seg_16_5_local_g2_0_64820;
  assign net_64822 = seg_16_5_local_g2_2_64822;
  assign net_64823 = seg_16_5_local_g2_3_64823;
  assign net_64826 = seg_16_5_local_g2_6_64826;
  assign net_64829 = seg_16_5_local_g3_1_64829;
  assign net_64830 = seg_16_5_local_g3_2_64830;
  assign net_64834 = seg_16_5_local_g3_6_64834;
  assign net_64835 = seg_16_5_local_g3_7_64835;
  assign net_64929 = seg_16_6_local_g0_2_64929;
  assign net_64931 = seg_16_6_local_g0_4_64931;
  assign net_64932 = seg_16_6_local_g0_5_64932;
  assign net_64933 = seg_16_6_local_g0_6_64933;
  assign net_64938 = seg_16_6_local_g1_3_64938;
  assign net_64941 = seg_16_6_local_g1_6_64941;
  assign net_64946 = seg_16_6_local_g2_3_64946;
  assign net_64952 = seg_16_6_local_g3_1_64952;
  assign net_64956 = seg_16_6_local_g3_5_64956;
  assign net_65050 = seg_16_7_local_g0_0_65050;
  assign net_65052 = seg_16_7_local_g0_2_65052;
  assign net_65053 = seg_16_7_local_g0_3_65053;
  assign net_65054 = seg_16_7_local_g0_4_65054;
  assign net_65062 = seg_16_7_local_g1_4_65062;
  assign net_65065 = seg_16_7_local_g1_7_65065;
  assign net_65070 = seg_16_7_local_g2_4_65070;
  assign net_65073 = seg_16_7_local_g2_7_65073;
  assign net_65176 = seg_16_8_local_g0_3_65176;
  assign net_65180 = seg_16_8_local_g0_7_65180;
  assign net_65185 = seg_16_8_local_g1_4_65185;
  assign net_65186 = seg_16_8_local_g1_5_65186;
  assign net_65303 = seg_16_9_local_g0_7_65303;
  assign net_65304 = seg_16_9_local_g1_0_65304;
  assign net_65307 = seg_16_9_local_g1_3_65307;
  assign net_65310 = seg_16_9_local_g1_6_65310;
  assign net_65319 = seg_16_9_local_g2_7_65319;
  assign net_65327 = seg_16_9_local_g3_7_65327;
  assign net_65421 = seg_16_10_local_g0_2_65421;
  assign net_65423 = seg_16_10_local_g0_4_65423;
  assign net_65427 = seg_16_10_local_g1_0_65427;
  assign net_65428 = seg_16_10_local_g1_1_65428;
  assign net_65436 = seg_16_10_local_g2_1_65436;
  assign net_65438 = seg_16_10_local_g2_3_65438;
  assign net_65439 = seg_16_10_local_g2_4_65439;
  assign net_65444 = seg_16_10_local_g3_1_65444;
  assign net_65445 = seg_16_10_local_g3_2_65445;
  assign net_65446 = seg_16_10_local_g3_3_65446;
  assign net_65543 = seg_16_11_local_g0_1_65543;
  assign net_65544 = seg_16_11_local_g0_2_65544;
  assign net_65546 = seg_16_11_local_g0_4_65546;
  assign net_65547 = seg_16_11_local_g0_5_65547;
  assign net_65555 = seg_16_11_local_g1_5_65555;
  assign net_65562 = seg_16_11_local_g2_4_65562;
  assign net_65565 = seg_16_11_local_g2_7_65565;
  assign net_65567 = seg_16_11_local_g3_1_65567;
  assign net_65568 = seg_16_11_local_g3_2_65568;
  assign net_65569 = seg_16_11_local_g3_3_65569;
  assign net_65571 = seg_16_11_local_g3_5_65571;
  assign net_65572 = seg_16_11_local_g3_6_65572;
  assign net_65573 = seg_16_11_local_g3_7_65573;
  assign net_65667 = seg_16_12_local_g0_2_65667;
  assign net_65668 = seg_16_12_local_g0_3_65668;
  assign net_65670 = seg_16_12_local_g0_5_65670;
  assign net_65672 = seg_16_12_local_g0_7_65672;
  assign net_65673 = seg_16_12_local_g1_0_65673;
  assign net_65674 = seg_16_12_local_g1_1_65674;
  assign net_65677 = seg_16_12_local_g1_4_65677;
  assign net_65678 = seg_16_12_local_g1_5_65678;
  assign net_65679 = seg_16_12_local_g1_6_65679;
  assign net_65680 = seg_16_12_local_g1_7_65680;
  assign net_65682 = seg_16_12_local_g2_1_65682;
  assign net_65686 = seg_16_12_local_g2_5_65686;
  assign net_65690 = seg_16_12_local_g3_1_65690;
  assign net_65694 = seg_16_12_local_g3_5_65694;
  assign net_65790 = seg_16_13_local_g0_2_65790;
  assign net_65792 = seg_16_13_local_g0_4_65792;
  assign net_65796 = seg_16_13_local_g1_0_65796;
  assign net_65797 = seg_16_13_local_g1_1_65797;
  assign net_65799 = seg_16_13_local_g1_3_65799;
  assign net_65800 = seg_16_13_local_g1_4_65800;
  assign net_65806 = seg_16_13_local_g2_2_65806;
  assign net_65807 = seg_16_13_local_g2_3_65807;
  assign net_65810 = seg_16_13_local_g2_6_65810;
  assign net_65812 = seg_16_13_local_g3_0_65812;
  assign net_65813 = seg_16_13_local_g3_1_65813;
  assign net_65814 = seg_16_13_local_g3_2_65814;
  assign net_65815 = seg_16_13_local_g3_3_65815;
  assign net_65816 = seg_16_13_local_g3_4_65816;
  assign net_65819 = seg_16_13_local_g3_7_65819;
  assign net_65911 = seg_16_14_local_g0_0_65911;
  assign net_65912 = seg_16_14_local_g0_1_65912;
  assign net_65913 = seg_16_14_local_g0_2_65913;
  assign net_65917 = seg_16_14_local_g0_6_65917;
  assign net_65919 = seg_16_14_local_g1_0_65919;
  assign net_65923 = seg_16_14_local_g1_4_65923;
  assign net_65924 = seg_16_14_local_g1_5_65924;
  assign net_65925 = seg_16_14_local_g1_6_65925;
  assign net_65926 = seg_16_14_local_g1_7_65926;
  assign net_65930 = seg_16_14_local_g2_3_65930;
  assign net_65933 = seg_16_14_local_g2_6_65933;
  assign net_65934 = seg_16_14_local_g2_7_65934;
  assign net_65935 = seg_16_14_local_g3_0_65935;
  assign net_65937 = seg_16_14_local_g3_2_65937;
  assign net_65938 = seg_16_14_local_g3_3_65938;
  assign net_65940 = seg_16_14_local_g3_5_65940;
  assign net_66040 = seg_16_15_local_g0_6_66040;
  assign net_66041 = seg_16_15_local_g0_7_66041;
  assign net_66049 = seg_16_15_local_g1_7_66049;
  assign net_66050 = seg_16_15_local_g2_0_66050;
  assign net_66051 = seg_16_15_local_g2_1_66051;
  assign net_66054 = seg_16_15_local_g2_4_66054;
  assign net_66063 = seg_16_15_local_g3_5_66063;
  assign net_66064 = seg_16_15_local_g3_6_66064;
  assign net_66160 = seg_16_16_local_g0_3_66160;
  assign net_66161 = seg_16_16_local_g0_4_66161;
  assign net_66162 = seg_16_16_local_g0_5_66162;
  assign net_66164 = seg_16_16_local_g0_7_66164;
  assign net_66165 = seg_16_16_local_g1_0_66165;
  assign net_66167 = seg_16_16_local_g1_2_66167;
  assign net_66169 = seg_16_16_local_g1_4_66169;
  assign net_66171 = seg_16_16_local_g1_6_66171;
  assign net_66172 = seg_16_16_local_g1_7_66172;
  assign net_66176 = seg_16_16_local_g2_3_66176;
  assign net_66180 = seg_16_16_local_g2_7_66180;
  assign net_66185 = seg_16_16_local_g3_4_66185;
  assign net_66187 = seg_16_16_local_g3_6_66187;
  assign net_66188 = seg_16_16_local_g3_7_66188;
  assign net_66280 = seg_16_17_local_g0_0_66280;
  assign net_66282 = seg_16_17_local_g0_2_66282;
  assign net_66283 = seg_16_17_local_g0_3_66283;
  assign net_66284 = seg_16_17_local_g0_4_66284;
  assign net_66293 = seg_16_17_local_g1_5_66293;
  assign net_66297 = seg_16_17_local_g2_1_66297;
  assign net_66299 = seg_16_17_local_g2_3_66299;
  assign net_66302 = seg_16_17_local_g2_6_66302;
  assign net_66303 = seg_16_17_local_g2_7_66303;
  assign net_66304 = seg_16_17_local_g3_0_66304;
  assign net_66305 = seg_16_17_local_g3_1_66305;
  assign net_66308 = seg_16_17_local_g3_4_66308;
  assign net_66310 = seg_16_17_local_g3_6_66310;
  assign net_66414 = seg_16_18_local_g1_3_66414;
  assign net_66425 = seg_16_18_local_g2_6_66425;
  assign net_6717 = seg_1_1_local_g0_2_6717;
  assign net_6720 = seg_1_1_local_g0_5_6720;
  assign net_6721 = seg_1_1_local_g0_6_6721;
  assign net_6726 = seg_1_1_local_g1_3_6726;
  assign net_6727 = seg_1_1_local_g1_4_6727;
  assign net_6730 = seg_1_1_local_g1_7_6730;
  assign net_6745 = seg_1_1_local_g3_6_6745;
  assign net_68021 = seg_16_31_local_g0_6_68021;
  assign net_68025 = seg_16_31_local_g1_2_68025;
  assign net_68281 = seg_17_2_local_g1_7_68281;
  assign net_68292 = seg_17_2_local_g3_2_68292;
  assign net_68391 = seg_17_3_local_g0_2_68391;
  assign net_68392 = seg_17_3_local_g0_3_68392;
  assign net_68400 = seg_17_3_local_g1_3_68400;
  assign net_68409 = seg_17_3_local_g2_4_68409;
  assign net_68413 = seg_17_3_local_g3_0_68413;
  assign net_68515 = seg_17_4_local_g0_3_68515;
  assign net_68520 = seg_17_4_local_g1_0_68520;
  assign net_68522 = seg_17_4_local_g1_2_68522;
  assign net_68523 = seg_17_4_local_g1_3_68523;
  assign net_68525 = seg_17_4_local_g1_5_68525;
  assign net_68526 = seg_17_4_local_g1_6_68526;
  assign net_68527 = seg_17_4_local_g1_7_68527;
  assign net_68535 = seg_17_4_local_g2_7_68535;
  assign net_68638 = seg_17_5_local_g0_3_68638;
  assign net_68642 = seg_17_5_local_g0_7_68642;
  assign net_68643 = seg_17_5_local_g1_0_68643;
  assign net_68644 = seg_17_5_local_g1_1_68644;
  assign net_68646 = seg_17_5_local_g1_3_68646;
  assign net_68653 = seg_17_5_local_g2_2_68653;
  assign net_68666 = seg_17_5_local_g3_7_68666;
  assign net_68764 = seg_17_6_local_g0_6_68764;
  assign net_68771 = seg_17_6_local_g1_5_68771;
  assign net_68779 = seg_17_6_local_g2_5_68779;
  assign net_68783 = seg_17_6_local_g3_1_68783;
  assign net_68785 = seg_17_6_local_g3_3_68785;
  assign net_68888 = seg_17_7_local_g0_7_68888;
  assign net_68899 = seg_17_7_local_g2_2_68899;
  assign net_69005 = seg_17_8_local_g0_1_69005;
  assign net_69006 = seg_17_8_local_g0_2_69006;
  assign net_69009 = seg_17_8_local_g0_5_69009;
  assign net_69013 = seg_17_8_local_g1_1_69013;
  assign net_69014 = seg_17_8_local_g1_2_69014;
  assign net_69019 = seg_17_8_local_g1_7_69019;
  assign net_69020 = seg_17_8_local_g2_0_69020;
  assign net_69022 = seg_17_8_local_g2_2_69022;
  assign net_69024 = seg_17_8_local_g2_4_69024;
  assign net_69028 = seg_17_8_local_g3_0_69028;
  assign net_69030 = seg_17_8_local_g3_2_69030;
  assign net_69032 = seg_17_8_local_g3_4_69032;
  assign net_6904 = seg_1_2_local_g0_2_6904;
  assign net_6905 = seg_1_2_local_g0_3_6905;
  assign net_6907 = seg_1_2_local_g0_5_6907;
  assign net_6909 = seg_1_2_local_g0_7_6909;
  assign net_6912 = seg_1_2_local_g1_2_6912;
  assign net_69128 = seg_17_9_local_g0_1_69128;
  assign net_69131 = seg_17_9_local_g0_4_69131;
  assign net_6915 = seg_1_2_local_g1_5_6915;
  assign net_6917 = seg_1_2_local_g1_7_6917;
  assign net_6919 = seg_1_2_local_g2_1_6919;
  assign net_6922 = seg_1_2_local_g2_4_6922;
  assign net_6924 = seg_1_2_local_g2_6_6924;
  assign net_6925 = seg_1_2_local_g2_7_6925;
  assign net_69254 = seg_17_10_local_g0_4_69254;
  assign net_69258 = seg_17_10_local_g1_0_69258;
  assign net_69263 = seg_17_10_local_g1_5_69263;
  assign net_69265 = seg_17_10_local_g1_7_69265;
  assign net_69269 = seg_17_10_local_g2_3_69269;
  assign net_69270 = seg_17_10_local_g2_4_69270;
  assign net_69280 = seg_17_10_local_g3_6_69280;
  assign net_69373 = seg_17_11_local_g0_0_69373;
  assign net_69374 = seg_17_11_local_g0_1_69374;
  assign net_69378 = seg_17_11_local_g0_5_69378;
  assign net_69380 = seg_17_11_local_g0_7_69380;
  assign net_69381 = seg_17_11_local_g1_0_69381;
  assign net_69384 = seg_17_11_local_g1_3_69384;
  assign net_69385 = seg_17_11_local_g1_4_69385;
  assign net_69386 = seg_17_11_local_g1_5_69386;
  assign net_69388 = seg_17_11_local_g1_7_69388;
  assign net_69389 = seg_17_11_local_g2_0_69389;
  assign net_69391 = seg_17_11_local_g2_2_69391;
  assign net_69395 = seg_17_11_local_g2_6_69395;
  assign net_69397 = seg_17_11_local_g3_0_69397;
  assign net_69399 = seg_17_11_local_g3_2_69399;
  assign net_69402 = seg_17_11_local_g3_5_69402;
  assign net_69403 = seg_17_11_local_g3_6_69403;
  assign net_69499 = seg_17_12_local_g0_3_69499;
  assign net_69509 = seg_17_12_local_g1_5_69509;
  assign net_69515 = seg_17_12_local_g2_3_69515;
  assign net_69518 = seg_17_12_local_g2_6_69518;
  assign net_69521 = seg_17_12_local_g3_1_69521;
  assign net_69522 = seg_17_12_local_g3_2_69522;
  assign net_69525 = seg_17_12_local_g3_5_69525;
  assign net_69526 = seg_17_12_local_g3_6_69526;
  assign net_69623 = seg_17_13_local_g0_4_69623;
  assign net_69637 = seg_17_13_local_g2_2_69637;
  assign net_69638 = seg_17_13_local_g2_3_69638;
  assign net_69639 = seg_17_13_local_g2_4_69639;
  assign net_69641 = seg_17_13_local_g2_6_69641;
  assign net_69644 = seg_17_13_local_g3_1_69644;
  assign net_69646 = seg_17_13_local_g3_3_69646;
  assign net_69648 = seg_17_13_local_g3_5_69648;
  assign net_69650 = seg_17_13_local_g3_7_69650;
  assign net_69744 = seg_17_14_local_g0_2_69744;
  assign net_69746 = seg_17_14_local_g0_4_69746;
  assign net_69747 = seg_17_14_local_g0_5_69747;
  assign net_69748 = seg_17_14_local_g0_6_69748;
  assign net_69753 = seg_17_14_local_g1_3_69753;
  assign net_69754 = seg_17_14_local_g1_4_69754;
  assign net_69755 = seg_17_14_local_g1_5_69755;
  assign net_69756 = seg_17_14_local_g1_6_69756;
  assign net_69757 = seg_17_14_local_g1_7_69757;
  assign net_69758 = seg_17_14_local_g2_0_69758;
  assign net_69760 = seg_17_14_local_g2_2_69760;
  assign net_69762 = seg_17_14_local_g2_4_69762;
  assign net_69763 = seg_17_14_local_g2_5_69763;
  assign net_69764 = seg_17_14_local_g2_6_69764;
  assign net_69765 = seg_17_14_local_g2_7_69765;
  assign net_69766 = seg_17_14_local_g3_0_69766;
  assign net_69768 = seg_17_14_local_g3_2_69768;
  assign net_69770 = seg_17_14_local_g3_4_69770;
  assign net_69772 = seg_17_14_local_g3_6_69772;
  assign net_69773 = seg_17_14_local_g3_7_69773;
  assign net_69868 = seg_17_15_local_g0_3_69868;
  assign net_69882 = seg_17_15_local_g2_1_69882;
  assign net_69883 = seg_17_15_local_g2_2_69883;
  assign net_69884 = seg_17_15_local_g2_3_69884;
  assign net_69886 = seg_17_15_local_g2_5_69886;
  assign net_69891 = seg_17_15_local_g3_2_69891;
  assign net_69892 = seg_17_15_local_g3_3_69892;
  assign net_69894 = seg_17_15_local_g3_5_69894;
  assign net_69990 = seg_17_16_local_g0_2_69990;
  assign net_69991 = seg_17_16_local_g0_3_69991;
  assign net_69997 = seg_17_16_local_g1_1_69997;
  assign net_70000 = seg_17_16_local_g1_4_70000;
  assign net_70001 = seg_17_16_local_g1_5_70001;
  assign net_70002 = seg_17_16_local_g1_6_70002;
  assign net_70003 = seg_17_16_local_g1_7_70003;
  assign net_70008 = seg_17_16_local_g2_4_70008;
  assign net_70016 = seg_17_16_local_g3_4_70016;
  assign net_70111 = seg_17_17_local_g0_0_70111;
  assign net_70114 = seg_17_17_local_g0_3_70114;
  assign net_70115 = seg_17_17_local_g0_4_70115;
  assign net_70116 = seg_17_17_local_g0_5_70116;
  assign net_70117 = seg_17_17_local_g0_6_70117;
  assign net_70118 = seg_17_17_local_g0_7_70118;
  assign net_70119 = seg_17_17_local_g1_0_70119;
  assign net_70120 = seg_17_17_local_g1_1_70120;
  assign net_70124 = seg_17_17_local_g1_5_70124;
  assign net_70131 = seg_17_17_local_g2_4_70131;
  assign net_70134 = seg_17_17_local_g2_7_70134;
  assign net_70138 = seg_17_17_local_g3_3_70138;
  assign net_70238 = seg_17_18_local_g0_4_70238;
  assign net_7050 = seg_1_3_local_g0_1_7050;
  assign net_7052 = seg_1_3_local_g0_3_7052;
  assign net_7056 = seg_1_3_local_g0_7_7056;
  assign net_7057 = seg_1_3_local_g1_0_7057;
  assign net_7058 = seg_1_3_local_g1_1_7058;
  assign net_7060 = seg_1_3_local_g1_3_7060;
  assign net_7062 = seg_1_3_local_g1_5_7062;
  assign net_7065 = seg_1_3_local_g2_0_7065;
  assign net_7066 = seg_1_3_local_g2_1_7066;
  assign net_7072 = seg_1_3_local_g2_7_7072;
  assign net_7074 = seg_1_3_local_g3_1_7074;
  assign net_7075 = seg_1_3_local_g3_2_7075;
  assign net_7077 = seg_1_3_local_g3_4_7077;
  assign net_7078 = seg_1_3_local_g3_5_7078;
  assign net_71855 = seg_17_31_local_g1_1_71855;
  assign net_71884 = seg_18_0_local_g1_0_71884;
  assign net_7196 = seg_1_4_local_g0_0_7196;
  assign net_7199 = seg_1_4_local_g0_3_7199;
  assign net_7201 = seg_1_4_local_g0_5_7201;
  assign net_7205 = seg_1_4_local_g1_1_7205;
  assign net_7207 = seg_1_4_local_g1_3_7207;
  assign net_7209 = seg_1_4_local_g1_5_7209;
  assign net_72103 = seg_18_2_local_g0_6_72103;
  assign net_72109 = seg_18_2_local_g1_4_72109;
  assign net_72116 = seg_18_2_local_g2_3_72116;
  assign net_7213 = seg_1_4_local_g2_1_7213;
  assign net_7214 = seg_1_4_local_g2_2_7214;
  assign net_7218 = seg_1_4_local_g2_6_7218;
  assign net_7222 = seg_1_4_local_g3_2_7222;
  assign net_72222 = seg_18_3_local_g0_2_72222;
  assign net_72223 = seg_18_3_local_g0_3_72223;
  assign net_72224 = seg_18_3_local_g0_4_72224;
  assign net_72228 = seg_18_3_local_g1_0_72228;
  assign net_72229 = seg_18_3_local_g1_1_72229;
  assign net_72233 = seg_18_3_local_g1_5_72233;
  assign net_72235 = seg_18_3_local_g1_7_72235;
  assign net_72249 = seg_18_3_local_g3_5_72249;
  assign net_7226 = seg_1_4_local_g3_6_7226;
  assign net_72344 = seg_18_4_local_g0_1_72344;
  assign net_72345 = seg_18_4_local_g0_2_72345;
  assign net_72346 = seg_18_4_local_g0_3_72346;
  assign net_72347 = seg_18_4_local_g0_4_72347;
  assign net_72349 = seg_18_4_local_g0_6_72349;
  assign net_72350 = seg_18_4_local_g0_7_72350;
  assign net_72351 = seg_18_4_local_g1_0_72351;
  assign net_72352 = seg_18_4_local_g1_1_72352;
  assign net_72353 = seg_18_4_local_g1_2_72353;
  assign net_72354 = seg_18_4_local_g1_3_72354;
  assign net_72355 = seg_18_4_local_g1_4_72355;
  assign net_72356 = seg_18_4_local_g1_5_72356;
  assign net_72358 = seg_18_4_local_g1_7_72358;
  assign net_72359 = seg_18_4_local_g2_0_72359;
  assign net_72360 = seg_18_4_local_g2_1_72360;
  assign net_72364 = seg_18_4_local_g2_5_72364;
  assign net_72469 = seg_18_5_local_g0_3_72469;
  assign net_72470 = seg_18_5_local_g0_4_72470;
  assign net_72472 = seg_18_5_local_g0_6_72472;
  assign net_72474 = seg_18_5_local_g1_0_72474;
  assign net_72475 = seg_18_5_local_g1_1_72475;
  assign net_72477 = seg_18_5_local_g1_3_72477;
  assign net_72478 = seg_18_5_local_g1_4_72478;
  assign net_72479 = seg_18_5_local_g1_5_72479;
  assign net_72482 = seg_18_5_local_g2_0_72482;
  assign net_72495 = seg_18_5_local_g3_5_72495;
  assign net_72590 = seg_18_6_local_g0_1_72590;
  assign net_72594 = seg_18_6_local_g0_5_72594;
  assign net_72597 = seg_18_6_local_g1_0_72597;
  assign net_72598 = seg_18_6_local_g1_1_72598;
  assign net_72599 = seg_18_6_local_g1_2_72599;
  assign net_72604 = seg_18_6_local_g1_7_72604;
  assign net_72612 = seg_18_6_local_g2_7_72612;
  assign net_72618 = seg_18_6_local_g3_5_72618;
  assign net_72717 = seg_18_7_local_g0_5_72717;
  assign net_72718 = seg_18_7_local_g0_6_72718;
  assign net_72719 = seg_18_7_local_g0_7_72719;
  assign net_72721 = seg_18_7_local_g1_1_72721;
  assign net_72723 = seg_18_7_local_g1_3_72723;
  assign net_72725 = seg_18_7_local_g1_5_72725;
  assign net_72727 = seg_18_7_local_g1_7_72727;
  assign net_72728 = seg_18_7_local_g2_0_72728;
  assign net_72730 = seg_18_7_local_g2_2_72730;
  assign net_72734 = seg_18_7_local_g2_6_72734;
  assign net_72742 = seg_18_7_local_g3_6_72742;
  assign net_72836 = seg_18_8_local_g0_1_72836;
  assign net_72840 = seg_18_8_local_g0_5_72840;
  assign net_72846 = seg_18_8_local_g1_3_72846;
  assign net_72848 = seg_18_8_local_g1_5_72848;
  assign net_72850 = seg_18_8_local_g1_7_72850;
  assign net_72854 = seg_18_8_local_g2_3_72854;
  assign net_72970 = seg_18_9_local_g1_4_72970;
  assign net_72971 = seg_18_9_local_g1_5_72971;
  assign net_72973 = seg_18_9_local_g1_7_72973;
  assign net_72974 = seg_18_9_local_g2_0_72974;
  assign net_72976 = seg_18_9_local_g2_2_72976;
  assign net_72987 = seg_18_9_local_g3_5_72987;
  assign net_73081 = seg_18_10_local_g0_0_73081;
  assign net_73082 = seg_18_10_local_g0_1_73082;
  assign net_73086 = seg_18_10_local_g0_5_73086;
  assign net_73087 = seg_18_10_local_g0_6_73087;
  assign net_73091 = seg_18_10_local_g1_2_73091;
  assign net_73094 = seg_18_10_local_g1_5_73094;
  assign net_73095 = seg_18_10_local_g1_6_73095;
  assign net_73096 = seg_18_10_local_g1_7_73096;
  assign net_73097 = seg_18_10_local_g2_0_73097;
  assign net_73103 = seg_18_10_local_g2_6_73103;
  assign net_73104 = seg_18_10_local_g2_7_73104;
  assign net_73106 = seg_18_10_local_g3_1_73106;
  assign net_73107 = seg_18_10_local_g3_2_73107;
  assign net_73205 = seg_18_11_local_g0_1_73205;
  assign net_73210 = seg_18_11_local_g0_6_73210;
  assign net_73211 = seg_18_11_local_g0_7_73211;
  assign net_73218 = seg_18_11_local_g1_6_73218;
  assign net_73220 = seg_18_11_local_g2_0_73220;
  assign net_73223 = seg_18_11_local_g2_3_73223;
  assign net_73225 = seg_18_11_local_g2_5_73225;
  assign net_73228 = seg_18_11_local_g3_0_73228;
  assign net_73330 = seg_18_12_local_g0_3_73330;
  assign net_73331 = seg_18_12_local_g0_4_73331;
  assign net_73335 = seg_18_12_local_g1_0_73335;
  assign net_73336 = seg_18_12_local_g1_1_73336;
  assign net_73342 = seg_18_12_local_g1_7_73342;
  assign net_73352 = seg_18_12_local_g3_1_73352;
  assign net_73353 = seg_18_12_local_g3_2_73353;
  assign net_7343 = seg_1_5_local_g0_0_7343;
  assign net_73451 = seg_18_13_local_g0_1_73451;
  assign net_73459 = seg_18_13_local_g1_1_73459;
  assign net_7346 = seg_1_5_local_g0_3_7346;
  assign net_73467 = seg_18_13_local_g2_1_73467;
  assign net_73475 = seg_18_13_local_g3_1_73475;
  assign net_73477 = seg_18_13_local_g3_3_73477;
  assign net_73481 = seg_18_13_local_g3_7_73481;
  assign net_7349 = seg_1_5_local_g0_6_7349;
  assign net_7353 = seg_1_5_local_g1_2_7353;
  assign net_7357 = seg_1_5_local_g1_6_7357;
  assign net_73573 = seg_18_14_local_g0_0_73573;
  assign net_73575 = seg_18_14_local_g0_2_73575;
  assign net_73576 = seg_18_14_local_g0_3_73576;
  assign net_73582 = seg_18_14_local_g1_1_73582;
  assign net_73584 = seg_18_14_local_g1_3_73584;
  assign net_73587 = seg_18_14_local_g1_6_73587;
  assign net_7359 = seg_1_5_local_g2_0_7359;
  assign net_73590 = seg_18_14_local_g2_1_73590;
  assign net_73599 = seg_18_14_local_g3_2_73599;
  assign net_7361 = seg_1_5_local_g2_2_7361;
  assign net_7363 = seg_1_5_local_g2_4_7363;
  assign net_7364 = seg_1_5_local_g2_5_7364;
  assign net_7366 = seg_1_5_local_g2_7_7366;
  assign net_73697 = seg_18_15_local_g0_1_73697;
  assign net_73698 = seg_18_15_local_g0_2_73698;
  assign net_73700 = seg_18_15_local_g0_4_73700;
  assign net_73701 = seg_18_15_local_g0_5_73701;
  assign net_73702 = seg_18_15_local_g0_6_73702;
  assign net_73703 = seg_18_15_local_g0_7_73703;
  assign net_73704 = seg_18_15_local_g1_0_73704;
  assign net_73705 = seg_18_15_local_g1_1_73705;
  assign net_73706 = seg_18_15_local_g1_2_73706;
  assign net_73707 = seg_18_15_local_g1_3_73707;
  assign net_73708 = seg_18_15_local_g1_4_73708;
  assign net_73709 = seg_18_15_local_g1_5_73709;
  assign net_73711 = seg_18_15_local_g1_7_73711;
  assign net_73722 = seg_18_15_local_g3_2_73722;
  assign net_73723 = seg_18_15_local_g3_3_73723;
  assign net_73724 = seg_18_15_local_g3_4_73724;
  assign net_73819 = seg_18_16_local_g0_0_73819;
  assign net_73830 = seg_18_16_local_g1_3_73830;
  assign net_73835 = seg_18_16_local_g2_0_73835;
  assign net_73839 = seg_18_16_local_g2_4_73839;
  assign net_73841 = seg_18_16_local_g2_6_73841;
  assign net_73843 = seg_18_16_local_g3_0_73843;
  assign net_73844 = seg_18_16_local_g3_1_73844;
  assign net_73848 = seg_18_16_local_g3_5_73848;
  assign net_73850 = seg_18_16_local_g3_7_73850;
  assign net_73973 = seg_18_17_local_g3_7_73973;
  assign net_7491 = seg_1_6_local_g0_1_7491;
  assign net_7506 = seg_1_6_local_g2_0_7506;
  assign net_7509 = seg_1_6_local_g2_3_7509;
  assign net_7510 = seg_1_6_local_g2_4_7510;
  assign net_7519 = seg_1_6_local_g3_5_7519;
  assign net_75679 = seg_18_31_local_g0_2_75679;
  assign net_75682 = seg_18_31_local_g0_5_75682;
  assign net_7648 = seg_1_7_local_g1_3_7648;
  assign net_7651 = seg_1_7_local_g1_6_7651;
  assign net_7792 = seg_1_8_local_g1_0_7792;
  assign net_7798 = seg_1_8_local_g1_6_7798;
  assign net_7801 = seg_1_8_local_g2_1_7801;
  assign net_7802 = seg_1_8_local_g2_2_7802;
  assign net_7806 = seg_1_8_local_g2_6_7806;
  assign net_7808 = seg_1_8_local_g3_0_7808;
  assign net_7812 = seg_1_8_local_g3_4_7812;
  assign net_7815 = seg_1_8_local_g3_7_7815;
  assign net_79130 = seg_20_2_local_g0_2_79130;
  assign net_79143 = seg_20_2_local_g1_7_79143;
  assign net_79155 = seg_20_2_local_g3_3_79155;
  assign net_79259 = seg_20_3_local_g1_0_79259;
  assign net_79260 = seg_20_3_local_g1_1_79260;
  assign net_79268 = seg_20_3_local_g2_1_79268;
  assign net_79270 = seg_20_3_local_g2_3_79270;
  assign net_79278 = seg_20_3_local_g3_3_79278;
  assign net_79279 = seg_20_3_local_g3_4_79279;
  assign net_7931 = seg_1_9_local_g0_0_7931;
  assign net_7936 = seg_1_9_local_g0_5_7936;
  assign net_79387 = seg_20_4_local_g1_5_79387;
  assign net_79388 = seg_20_4_local_g1_6_79388;
  assign net_79401 = seg_20_4_local_g3_3_79401;
  assign net_7944 = seg_1_9_local_g1_5_7944;
  assign net_7946 = seg_1_9_local_g1_7_7946;
  assign net_79501 = seg_20_5_local_g0_4_79501;
  assign net_79504 = seg_20_5_local_g0_7_79504;
  assign net_79505 = seg_20_5_local_g1_0_79505;
  assign net_79508 = seg_20_5_local_g1_3_79508;
  assign net_79519 = seg_20_5_local_g2_6_79519;
  assign net_79522 = seg_20_5_local_g3_1_79522;
  assign net_79527 = seg_20_5_local_g3_6_79527;
  assign net_79528 = seg_20_5_local_g3_7_79528;
  assign net_7956 = seg_1_9_local_g3_1_7956;
  assign net_7960 = seg_1_9_local_g3_5_7960;
  assign net_7961 = seg_1_9_local_g3_6_7961;
  assign net_7962 = seg_1_9_local_g3_7_7962;
  assign net_79630 = seg_20_6_local_g1_2_79630;
  assign net_79631 = seg_20_6_local_g1_3_79631;
  assign net_79632 = seg_20_6_local_g1_4_79632;
  assign net_79633 = seg_20_6_local_g1_5_79633;
  assign net_79640 = seg_20_6_local_g2_4_79640;
  assign net_79641 = seg_20_6_local_g2_5_79641;
  assign net_79642 = seg_20_6_local_g2_6_79642;
  assign net_79645 = seg_20_6_local_g3_1_79645;
  assign net_79646 = seg_20_6_local_g3_2_79646;
  assign net_79647 = seg_20_6_local_g3_3_79647;
  assign net_79649 = seg_20_6_local_g3_5_79649;
  assign net_79745 = seg_20_7_local_g0_2_79745;
  assign net_79750 = seg_20_7_local_g0_7_79750;
  assign net_79752 = seg_20_7_local_g1_1_79752;
  assign net_79757 = seg_20_7_local_g1_6_79757;
  assign net_79770 = seg_20_7_local_g3_3_79770;
  assign net_79893 = seg_20_8_local_g3_3_79893;
  assign net_79996 = seg_20_9_local_g0_7_79996;
  assign net_79998 = seg_20_9_local_g1_1_79998;
  assign net_8 = seg_14_4_glb_netwk_3_8;
  assign net_80004 = seg_20_9_local_g1_7_80004;
  assign net_80020 = seg_20_9_local_g3_7_80020;
  assign net_80113 = seg_20_10_local_g0_1_80113;
  assign net_80114 = seg_20_10_local_g0_2_80114;
  assign net_80118 = seg_20_10_local_g0_6_80118;
  assign net_80119 = seg_20_10_local_g0_7_80119;
  assign net_80126 = seg_20_10_local_g1_6_80126;
  assign net_80127 = seg_20_10_local_g1_7_80127;
  assign net_80242 = seg_20_11_local_g0_7_80242;
  assign net_80244 = seg_20_11_local_g1_1_80244;
  assign net_80362 = seg_20_12_local_g0_4_80362;
  assign net_80383 = seg_20_12_local_g3_1_80383;
  assign net_80615 = seg_20_14_local_g1_3_80615;
  assign net_80631 = seg_20_14_local_g3_3_80631;
  assign net_8081 = seg_1_10_local_g0_3_8081;
  assign net_8083 = seg_1_10_local_g0_5_8083;
  assign net_8085 = seg_1_10_local_g0_7_8085;
  assign net_8089 = seg_1_10_local_g1_3_8089;
  assign net_8095 = seg_1_10_local_g2_1_8095;
  assign net_8098 = seg_1_10_local_g2_4_8098;
  assign net_8104 = seg_1_10_local_g3_2_8104;
  assign net_8108 = seg_1_10_local_g3_6_8108;
  assign net_8228 = seg_1_11_local_g0_3_8228;
  assign net_8232 = seg_1_11_local_g0_7_8232;
  assign net_8235 = seg_1_11_local_g1_2_8235;
  assign net_8246 = seg_1_11_local_g2_5_8246;
  assign net_8247 = seg_1_11_local_g2_6_8247;
  assign net_8248 = seg_1_11_local_g2_7_8248;
  assign net_8252 = seg_1_11_local_g3_3_8252;
  assign net_8254 = seg_1_11_local_g3_5_8254;
  assign net_82750 = seg_21_0_local_g1_4_82750;
  assign net_83100 = seg_21_3_local_g2_2_83100;
  assign net_83102 = seg_21_3_local_g2_4_83102;
  assign net_83106 = seg_21_3_local_g3_0_83106;
  assign net_83112 = seg_21_3_local_g3_6_83112;
  assign net_83206 = seg_21_4_local_g0_1_83206;
  assign net_83219 = seg_21_4_local_g1_6_83219;
  assign net_83227 = seg_21_4_local_g2_6_83227;
  assign net_83228 = seg_21_4_local_g2_7_83228;
  assign net_83236 = seg_21_4_local_g3_7_83236;
  assign net_83328 = seg_21_5_local_g0_0_83328;
  assign net_83356 = seg_21_5_local_g3_4_83356;
  assign net_83357 = seg_21_5_local_g3_5_83357;
  assign net_83452 = seg_21_6_local_g0_1_83452;
  assign net_83471 = seg_21_6_local_g2_4_83471;
  assign net_83479 = seg_21_6_local_g3_4_83479;
  assign net_83481 = seg_21_6_local_g3_6_83481;
  assign net_83576 = seg_21_7_local_g0_2_83576;
  assign net_83577 = seg_21_7_local_g0_3_83577;
  assign net_83579 = seg_21_7_local_g0_5_83579;
  assign net_83600 = seg_21_7_local_g3_2_83600;
  assign net_83699 = seg_21_8_local_g0_2_83699;
  assign net_83701 = seg_21_8_local_g0_4_83701;
  assign net_83703 = seg_21_8_local_g0_6_83703;
  assign net_83704 = seg_21_8_local_g0_7_83704;
  assign net_83706 = seg_21_8_local_g1_1_83706;
  assign net_83707 = seg_21_8_local_g1_2_83707;
  assign net_83710 = seg_21_8_local_g1_5_83710;
  assign net_83711 = seg_21_8_local_g1_6_83711;
  assign net_83716 = seg_21_8_local_g2_3_83716;
  assign net_83717 = seg_21_8_local_g2_4_83717;
  assign net_83719 = seg_21_8_local_g2_6_83719;
  assign net_83720 = seg_21_8_local_g2_7_83720;
  assign net_83721 = seg_21_8_local_g3_0_83721;
  assign net_83725 = seg_21_8_local_g3_4_83725;
  assign net_83726 = seg_21_8_local_g3_5_83726;
  assign net_83727 = seg_21_8_local_g3_6_83727;
  assign net_8375 = seg_1_12_local_g0_3_8375;
  assign net_8377 = seg_1_12_local_g0_5_8377;
  assign net_8378 = seg_1_12_local_g0_6_8378;
  assign net_8380 = seg_1_12_local_g1_0_8380;
  assign net_83825 = seg_21_9_local_g0_5_83825;
  assign net_8383 = seg_1_12_local_g1_3_8383;
  assign net_83830 = seg_21_9_local_g1_2_83830;
  assign net_83831 = seg_21_9_local_g1_3_83831;
  assign net_83832 = seg_21_9_local_g1_4_83832;
  assign net_83834 = seg_21_9_local_g1_6_83834;
  assign net_83835 = seg_21_9_local_g1_7_83835;
  assign net_83836 = seg_21_9_local_g2_0_83836;
  assign net_8384 = seg_1_12_local_g1_4_8384;
  assign net_83840 = seg_21_9_local_g2_4_83840;
  assign net_83847 = seg_21_9_local_g3_3_83847;
  assign net_83850 = seg_21_9_local_g3_6_83850;
  assign net_8392 = seg_1_12_local_g2_4_8392;
  assign net_83943 = seg_21_10_local_g0_0_83943;
  assign net_83951 = seg_21_10_local_g1_0_83951;
  assign net_83954 = seg_21_10_local_g1_3_83954;
  assign net_83956 = seg_21_10_local_g1_5_83956;
  assign net_83958 = seg_21_10_local_g1_7_83958;
  assign net_8519 = seg_1_13_local_g0_0_8519;
  assign net_8522 = seg_1_13_local_g0_3_8522;
  assign net_8525 = seg_1_13_local_g0_6_8525;
  assign net_8527 = seg_1_13_local_g1_0_8527;
  assign net_8529 = seg_1_13_local_g1_2_8529;
  assign net_8531 = seg_1_13_local_g1_4_8531;
  assign net_8533 = seg_1_13_local_g1_6_8533;
  assign net_8535 = seg_1_13_local_g2_0_8535;
  assign net_86583 = seg_22_0_local_g1_6_86583;
  assign net_8669 = seg_1_14_local_g0_3_8669;
  assign net_8670 = seg_1_14_local_g0_4_8670;
  assign net_8671 = seg_1_14_local_g0_5_8671;
  assign net_8673 = seg_1_14_local_g0_7_8673;
  assign net_8680 = seg_1_14_local_g1_6_8680;
  assign net_8683 = seg_1_14_local_g2_1_8683;
  assign net_8684 = seg_1_14_local_g2_2_8684;
  assign net_8689 = seg_1_14_local_g2_7_8689;
  assign net_86917 = seg_22_3_local_g0_4_86917;
  assign net_86924 = seg_22_3_local_g1_3_86924;
  assign net_86940 = seg_22_3_local_g3_3_86940;
  assign net_87036 = seg_22_4_local_g0_0_87036;
  assign net_87054 = seg_22_4_local_g2_2_87054;
  assign net_87059 = seg_22_4_local_g2_7_87059;
  assign net_87163 = seg_22_5_local_g0_4_87163;
  assign net_87176 = seg_22_5_local_g2_1_87176;
  assign net_87177 = seg_22_5_local_g2_2_87177;
  assign net_87178 = seg_22_5_local_g2_3_87178;
  assign net_87183 = seg_22_5_local_g3_0_87183;
  assign net_87301 = seg_22_6_local_g2_3_87301;
  assign net_87305 = seg_22_6_local_g2_7_87305;
  assign net_87413 = seg_22_7_local_g1_0_87413;
  assign net_87428 = seg_22_7_local_g2_7_87428;
  assign net_87430 = seg_22_7_local_g3_1_87430;
  assign net_87434 = seg_22_7_local_g3_5_87434;
  assign net_87539 = seg_22_8_local_g1_3_87539;
  assign net_87542 = seg_22_8_local_g1_6_87542;
  assign net_87543 = seg_22_8_local_g1_7_87543;
  assign net_87547 = seg_22_8_local_g2_3_87547;
  assign net_87550 = seg_22_8_local_g2_6_87550;
  assign net_87557 = seg_22_8_local_g3_5_87557;
  assign net_87665 = seg_22_9_local_g1_6_87665;
  assign net_87668 = seg_22_9_local_g2_1_87668;
  assign net_87676 = seg_22_9_local_g3_1_87676;
  assign net_87677 = seg_22_9_local_g3_2_87677;
  assign net_87682 = seg_22_9_local_g3_7_87682;
  assign net_8813 = seg_1_15_local_g0_0_8813;
  assign net_8824 = seg_1_15_local_g1_3_8824;
  assign net_8827 = seg_1_15_local_g1_6_8827;
  assign net_8829 = seg_1_15_local_g2_0_8829;
  assign net_8830 = seg_1_15_local_g2_1_8830;
  assign net_8835 = seg_1_15_local_g2_6_8835;
  assign net_8838 = seg_1_15_local_g3_1_8838;
  assign net_8841 = seg_1_15_local_g3_4_8841;
  assign net_8965 = seg_1_16_local_g0_5_8965;
  assign net_8977 = seg_1_16_local_g2_1_8977;
  assign net_8981 = seg_1_16_local_g2_5_8981;
  assign net_8982 = seg_1_16_local_g2_6_8982;
  assign net_8984 = seg_1_16_local_g3_0_8984;
  assign net_8988 = seg_1_16_local_g3_4_8988;
  assign net_8989 = seg_1_16_local_g3_5_8989;
  assign net_9 = seg_23_9_glb_netwk_4_9;
  assign net_90410 = seg_23_0_local_g1_2_90410;
  assign net_90991 = seg_23_5_local_g0_1_90991;
  assign net_91009 = seg_23_5_local_g2_3_91009;
  assign net_91014 = seg_23_5_local_g3_0_91014;
  assign net_91018 = seg_23_5_local_g3_4_91018;
  assign net_91021 = seg_23_5_local_g3_7_91021;
  assign net_9107 = seg_1_17_local_g0_0_9107;
  assign net_9108 = seg_1_17_local_g0_1_9108;
  assign net_9111 = seg_1_17_local_g0_4_9111;
  assign net_91133 = seg_23_6_local_g2_4_91133;
  assign net_91137 = seg_23_6_local_g3_0_91137;
  assign net_91141 = seg_23_6_local_g3_4_91141;
  assign net_9130 = seg_1_17_local_g2_7_9130;
  assign net_91380 = seg_23_8_local_g2_5_91380;
  assign net_91495 = seg_23_9_local_g1_5_91495;
  assign net_9256 = seg_1_18_local_g0_2_9256;
  assign net_9261 = seg_1_18_local_g0_7_9261;
  assign net_9267 = seg_1_18_local_g1_5_9267;
  assign net_9281 = seg_1_18_local_g3_3_9281;
  assign net_9402 = seg_1_19_local_g0_1_9402;
  assign net_9407 = seg_1_19_local_g0_6_9407;
  assign net_9416 = seg_1_19_local_g1_7_9416;
  assign net_9554 = seg_1_20_local_g0_6_9554;
  assign net_9560 = seg_1_20_local_g1_4_9560;
  assign net_9564 = seg_1_20_local_g2_0_9564;
  assign net_9576 = seg_1_20_local_g3_4_9576;
  assign net_9700 = seg_1_21_local_g0_5_9700;
  assign net_9721 = seg_1_21_local_g3_2_9721;
  assign net_9843 = seg_1_22_local_g0_1_9843;
  assign net_9848 = seg_1_22_local_g0_6_9848;
  assign net_9851 = seg_1_22_local_g1_1_9851;
  assign net_99370 = seg_25_6_local_g0_0_99370;
  assign net_99373 = seg_25_6_local_g0_3_99373;
  assign net_99380 = seg_25_6_local_g1_2_99380;
  assign net_99383 = seg_25_6_local_g1_5_99383;
  assign net_99385 = seg_25_6_local_g1_7_99385;
  assign net_99386 = seg_25_6_local_g2_0_99386;
  assign net_99388 = seg_25_6_local_g2_2_99388;
  assign net_99389 = seg_25_6_local_g2_3_99389;
  assign net_99391 = seg_25_6_local_g2_5_99391;
  assign net_99394 = seg_25_6_local_g3_0_99394;
  assign net_99395 = seg_25_6_local_g3_1_99395;
  assign net_99396 = seg_25_6_local_g3_2_99396;
  assign net_99398 = seg_25_6_local_g3_4_99398;
  assign net_99399 = seg_25_6_local_g3_5_99399;
  assign net_99400 = seg_25_6_local_g3_6_99400;
  assign net_99401 = seg_25_6_local_g3_7_99401;
  assign net_99520 = seg_25_7_local_g0_0_99520;
  assign net_99521 = seg_25_7_local_g0_1_99521;
  assign net_99523 = seg_25_7_local_g0_3_99523;
  assign net_99527 = seg_25_7_local_g0_7_99527;
  assign net_99529 = seg_25_7_local_g1_1_99529;
  assign net_99530 = seg_25_7_local_g1_2_99530;
  assign net_99532 = seg_25_7_local_g1_4_99532;
  assign net_99533 = seg_25_7_local_g1_5_99533;
  assign net_99534 = seg_25_7_local_g1_6_99534;
  assign net_99535 = seg_25_7_local_g1_7_99535;
  assign net_99536 = seg_25_7_local_g2_0_99536;
  assign net_99543 = seg_25_7_local_g2_7_99543;
  assign net_99544 = seg_25_7_local_g3_0_99544;
  assign net_99545 = seg_25_7_local_g3_1_99545;
  assign net_99547 = seg_25_7_local_g3_3_99547;
  assign net_99549 = seg_25_7_local_g3_5_99549;
  assign seg_0_10_sp12_h_r_0_2200 = seg_10_10_sp12_h_r_20_2200;
  assign seg_0_10_sp4_h_r_40_2273 = net_2273;
  assign seg_0_10_sp4_r_v_b_37_2287 = net_2287;
  assign seg_0_10_sp4_r_v_b_39_2289 = net_2289;
  assign seg_0_10_sp4_r_v_b_43_2293 = net_2293;
  assign seg_0_10_sp4_r_v_b_45_2295 = net_2295;
  assign seg_0_10_sp4_r_v_b_47_2297 = net_2297;
  assign seg_0_10_sp4_v_b_16_1656 = net_1656;
  assign seg_0_10_sp4_v_b_18_1658 = net_1658;
  assign seg_0_10_sp4_v_t_36_2298 = seg_0_13_sp4_v_b_12_2298;
  assign seg_0_10_sp4_v_t_47_2309 = seg_0_12_sp4_v_b_34_2309;
  assign seg_0_11_sp12_h_r_1_2407 = seg_11_11_sp12_h_r_22_2407;
  assign seg_0_11_sp4_h_r_0_2444 = net_2444;
  assign seg_0_11_sp4_h_r_10_2446 = net_2446;
  assign seg_0_11_sp4_h_r_12_2448 = net_2448;
  assign seg_0_11_sp4_h_r_2_2456 = net_2456;
  assign seg_0_11_sp4_h_r_46_2485 = net_2485;
  assign seg_0_11_sp4_h_r_4_2478 = net_2478;
  assign seg_0_11_sp4_h_r_6_2488 = net_2488;
  assign seg_0_11_sp4_h_r_7_2489 = seg_3_11_sp4_h_r_42_2489;
  assign seg_0_11_sp4_h_r_8_2490 = net_2490;
  assign seg_0_11_sp4_h_r_9_2491 = seg_3_11_sp4_h_r_44_2491;
  assign seg_0_11_sp4_r_v_b_0_1850 = seg_1_9_sp4_v_b_24_1850;
  assign seg_0_11_sp4_r_v_b_12_2076 = seg_1_9_sp4_v_b_36_2076;
  assign seg_0_11_sp4_r_v_b_8_1858 = seg_1_9_sp4_v_b_32_1858;
  assign seg_0_11_sp4_v_b_5_1656 = seg_0_10_sp4_v_b_16_1656;
  assign seg_0_11_sp4_v_b_7_1658 = seg_0_10_sp4_v_b_18_1658;
  assign seg_0_12_sp4_h_r_16_2660 = net_2660;
  assign seg_0_12_sp4_h_r_20_2665 = net_2665;
  assign seg_0_12_sp4_r_v_b_11_2086 = net_2086;
  assign seg_0_12_sp4_r_v_b_25_2492 = net_2492;
  assign seg_0_12_sp4_r_v_b_31_2498 = net_2498;
  assign seg_0_12_sp4_r_v_b_39_2703 = net_2703;
  assign seg_0_12_sp4_v_b_12_2088 = net_2088;
  assign seg_0_12_sp4_v_b_34_2309 = net_2309;
  assign seg_0_12_sp4_v_t_43_2719 = seg_0_16_sp4_v_b_6_2719;
  assign seg_0_12_sp4_v_t_45_2721 = seg_0_16_sp4_v_b_8_2721;
  assign seg_0_13_sp4_h_r_0_2861 = net_2861;
  assign seg_0_13_sp4_h_r_24_2878 = net_2878;
  assign seg_0_13_sp4_h_r_38_2893 = net_2893;
  assign seg_0_13_sp4_r_v_b_21_2501 = net_2501;
  assign seg_0_13_sp4_r_v_b_27_2702 = net_2702;
  assign seg_0_13_sp4_r_v_b_3_2288 = net_2288;
  assign seg_0_13_sp4_v_b_12_2298 = net_2298;
  assign seg_0_14_sp4_v_t_39_3151 = seg_0_16_sp4_v_b_26_3151;
  assign seg_0_14_sp4_v_t_45_3157 = seg_0_16_sp4_v_b_32_3157;
  assign seg_0_14_sp4_v_t_46_3158 = seg_0_17_sp4_v_b_22_3158;
  assign seg_0_15_sp4_h_r_10_3300 = net_3300;
  assign seg_0_15_sp4_h_r_14_3304 = net_3304;
  assign seg_0_15_sp4_h_r_16_3306 = net_3306;
  assign seg_0_15_sp4_h_r_18_3308 = net_3308;
  assign seg_0_15_sp4_h_r_8_3344 = net_3344;
  assign seg_0_15_sp4_r_v_b_23_2920 = net_2920;
  assign seg_0_15_sp4_v_b_20_2720 = net_2720;
  assign seg_0_15_sp4_v_b_28_2926 = net_2926;
  assign seg_0_15_sp4_v_t_40_3362 = seg_0_18_sp4_v_b_16_3362;
  assign seg_0_15_sp4_v_t_43_3365 = seg_0_17_sp4_v_b_30_3365;
  assign seg_0_16_sp4_h_r_18_3514 = net_3514;
  assign seg_0_16_sp4_r_v_b_13_3137 = net_3137;
  assign seg_0_16_sp4_r_v_b_15_3139 = net_3139;
  assign seg_0_16_sp4_r_v_b_5_2913 = net_2913;
  assign seg_0_16_sp4_v_b_26_3151 = net_3151;
  assign seg_0_16_sp4_v_b_32_3157 = net_3157;
  assign seg_0_16_sp4_v_b_6_2719 = net_2719;
  assign seg_0_16_sp4_v_b_8_2721 = net_2721;
  assign seg_0_16_sp4_v_b_9_2720 = seg_0_15_sp4_v_b_20_2720;
  assign seg_0_17_sp4_h_r_26_3731 = net_3731;
  assign seg_0_17_sp4_h_r_4_3746 = net_3746;
  assign seg_0_17_sp4_h_r_8_3758 = net_3758;
  assign seg_0_17_sp4_r_v_b_17_3351 = net_3351;
  assign seg_0_17_sp4_r_v_b_29_3556 = net_3556;
  assign seg_0_17_sp4_r_v_b_35_3562 = net_3562;
  assign seg_0_17_sp4_v_b_22_3158 = net_3158;
  assign seg_0_17_sp4_v_b_30_3365 = net_3365;
  assign seg_0_17_sp4_v_b_4_2926 = seg_0_15_sp4_v_b_28_2926;
  assign seg_0_18_sp4_h_r_6_3965 = net_3965;
  assign seg_0_18_sp4_r_v_b_11_3356 = net_3356;
  assign seg_0_18_sp4_r_v_b_13_3553 = net_3553;
  assign seg_0_18_sp4_r_v_b_19_3559 = net_3559;
  assign seg_0_18_sp4_r_v_b_5_3350 = net_3350;
  assign seg_0_18_sp4_r_v_b_9_3354 = net_3354;
  assign seg_0_18_sp4_v_b_16_3362 = net_3362;
  assign seg_0_20_sp4_v_t_36_4435 = seg_0_23_sp4_v_b_12_4435;
  assign seg_0_22_sp4_v_t_47_4900 = seg_0_26_sp4_v_b_10_4900;
  assign seg_0_23_sp4_h_r_0_5039 = net_5039;
  assign seg_0_23_sp4_r_v_b_11_4433 = net_4433;
  assign seg_0_23_sp4_r_v_b_15_4653 = net_4653;
  assign seg_0_23_sp4_r_v_b_3_4425 = net_4425;
  assign seg_0_23_sp4_r_v_b_5_4427 = net_4427;
  assign seg_0_23_sp4_r_v_b_7_4429 = net_4429;
  assign seg_0_23_sp4_r_v_b_9_4431 = net_4431;
  assign seg_0_23_sp4_v_b_12_4435 = net_4435;
  assign seg_0_24_sp4_h_r_22_5260 = net_5260;
  assign seg_0_24_sp4_r_v_b_11_4660 = net_4660;
  assign seg_0_24_sp4_r_v_b_15_4880 = net_4880;
  assign seg_0_24_sp4_r_v_b_1_4650 = net_4650;
  assign seg_0_24_sp4_r_v_b_29_5091 = net_5091;
  assign seg_0_24_sp4_r_v_b_35_5097 = net_5097;
  assign seg_0_24_sp4_r_v_b_5_4654 = net_4654;
  assign seg_0_24_sp4_r_v_b_9_4658 = net_4658;
  assign seg_0_25_sp4_h_r_0_5453 = net_5453;
  assign seg_0_25_sp4_h_r_26_5472 = net_5472;
  assign seg_0_25_sp4_h_r_6_5497 = net_5497;
  assign seg_0_25_sp4_h_r_8_5499 = net_5499;
  assign seg_0_25_sp4_r_v_b_13_5088 = net_5088;
  assign seg_0_25_sp4_r_v_b_31_5299 = net_5299;
  assign seg_0_25_sp4_r_v_b_3_4879 = net_4879;
  assign seg_0_25_sp4_r_v_b_5_4881 = net_4881;
  assign seg_0_26_sp4_h_r_28_5683 = net_5683;
  assign seg_0_26_sp4_r_v_b_17_5298 = net_5298;
  assign seg_0_26_sp4_r_v_b_21_5302 = net_5302;
  assign seg_0_26_sp4_r_v_b_35_5511 = net_5511;
  assign seg_0_26_sp4_r_v_b_7_5093 = net_5093;
  assign seg_0_26_sp4_r_v_b_9_5095 = net_5095;
  assign seg_0_26_sp4_v_b_10_4900 = net_4900;
  assign seg_0_4_sp4_v_t_39_1031 = seg_0_8_sp4_v_b_2_1031;
  assign seg_0_4_sp4_v_t_45_1037 = seg_0_8_sp4_v_b_8_1037;
  assign seg_0_5_sp4_h_r_0_1178 = net_1178;
  assign seg_0_5_sp4_h_r_11_1181 = seg_1_5_sp4_h_r_22_1181;
  assign seg_0_5_sp4_h_r_14_1184 = net_1184;
  assign seg_0_5_sp4_h_r_24_1195 = net_1195;
  assign seg_0_5_sp4_h_r_28_1199 = net_1199;
  assign seg_0_5_sp4_h_r_34_1206 = net_1206;
  assign seg_0_5_sp4_h_r_38_1210 = net_1210;
  assign seg_0_5_sp4_h_r_3_1201 = seg_1_5_sp4_h_r_14_1201;
  assign seg_0_5_sp4_h_r_7_1223 = seg_1_5_sp4_h_r_18_1223;
  assign seg_0_5_sp4_h_r_8_1224 = seg_2_5_sp4_h_r_32_1224;
  assign seg_0_5_sp4_r_v_b_21_798 = net_798;
  assign seg_0_5_sp4_v_b_26_804 = net_804;
  assign seg_0_6_sp4_h_r_0_1384 = net_1384;
  assign seg_0_6_sp4_h_r_44_1423 = net_1423;
  assign seg_0_6_sp4_h_r_4_1418 = net_1418;
  assign seg_0_6_sp4_h_r_8_1430 = net_1430;
  assign seg_0_6_sp4_r_v_b_15_1019 = net_1019;
  assign seg_0_6_sp4_r_v_b_19_1023 = net_1023;
  assign seg_0_6_sp4_r_v_b_27_1228 = net_1228;
  assign seg_0_6_sp4_v_b_22_811 = net_811;
  assign seg_0_6_sp4_v_t_39_1447 = seg_0_8_sp4_v_b_26_1447;
  assign seg_0_7_neigh_op_bnr_3_1133 = seg_1_6_lutff_3_out_1133;
  assign seg_0_7_neigh_op_bnr_6_1136 = seg_1_6_lutff_6_out_1136;
  assign seg_0_7_neigh_op_tnr_3_1547 = seg_1_8_lutff_3_out_1547;
  assign seg_0_7_neigh_op_tnr_4_1548 = seg_1_8_lutff_4_out_1548;
  assign seg_0_7_neigh_op_tnr_7_1551 = seg_1_8_lutff_7_out_1551;
  assign seg_0_7_sp12_h_r_1_1555 = seg_9_7_sp12_h_r_18_1555;
  assign seg_0_7_sp4_h_r_10_1594 = net_1594;
  assign seg_0_7_sp4_h_r_14_1598 = net_1598;
  assign seg_0_7_sp4_h_r_32_1618 = net_1618;
  assign seg_0_7_sp4_h_r_6_1636 = net_1636;
  assign seg_0_7_sp4_r_v_b_13_1227 = net_1227;
  assign seg_0_7_sp4_r_v_b_19_1233 = net_1233;
  assign seg_0_7_sp4_r_v_b_21_1235 = net_1235;
  assign seg_0_7_sp4_r_v_b_22_1236 = seg_1_5_sp4_v_b_46_1236;
  assign seg_0_7_sp4_r_v_b_41_1645 = net_1645;
  assign seg_0_7_sp4_v_b_11_811 = seg_0_6_sp4_v_b_22_811;
  assign seg_0_7_sp4_v_b_2_804 = seg_0_5_sp4_v_b_26_804;
  assign seg_0_8_sp12_h_r_1_1764 = seg_11_8_sp12_h_r_22_1764;
  assign seg_0_8_sp4_h_r_0_1801 = net_1801;
  assign seg_0_8_sp4_h_r_12_1805 = net_1805;
  assign seg_0_8_sp4_h_r_20_1814 = net_1814;
  assign seg_0_8_sp4_r_v_b_7_1232 = net_1232;
  assign seg_0_8_sp4_v_b_26_1447 = net_1447;
  assign seg_0_8_sp4_v_b_2_1031 = net_1031;
  assign seg_0_8_sp4_v_b_8_1037 = net_1037;
  assign seg_0_9_sp12_h_r_1_1991 = seg_5_9_sp12_h_r_10_1991;
  assign seg_0_9_sp4_h_r_5_2071 = seg_1_9_sp4_h_r_16_2071;
  assign seg_0_9_sp4_v_t_36_2088 = seg_0_12_sp4_v_b_12_2088;
  assign seg_10_10_lutff_1_out_38564 = net_38564;
  assign seg_10_10_lutff_3_out_38566 = net_38566;
  assign seg_10_10_lutff_5_out_38568 = net_38568;
  assign seg_10_10_sp12_h_r_1_42526 = seg_17_10_sp12_h_r_14_42526;
  assign seg_10_10_sp12_h_r_20_2200 = net_2200;
  assign seg_10_10_sp4_h_r_0_42529 = net_42529;
  assign seg_10_10_sp4_h_r_14_38703 = net_38703;
  assign seg_10_10_sp4_h_r_28_34873 = net_34873;
  assign seg_10_10_sp4_h_r_32_34877 = net_34877;
  assign seg_10_10_sp4_v_b_14_38466 = net_38466;
  assign seg_10_10_sp4_v_b_32_38596 = net_38596;
  assign seg_10_10_sp4_v_b_46_38720 = net_38720;
  assign seg_10_10_sp4_v_b_4_38346 = net_38346;
  assign seg_10_11_lutff_0_out_38686 = net_38686;
  assign seg_10_11_lutff_1_out_38687 = net_38687;
  assign seg_10_11_lutff_3_out_38689 = net_38689;
  assign seg_10_11_lutff_6_out_38692 = net_38692;
  assign seg_10_11_neigh_op_bnr_1_42395 = seg_11_10_lutff_1_out_42395;
  assign seg_10_11_neigh_op_bnr_7_42401 = seg_11_10_lutff_7_out_42401;
  assign seg_10_11_sp4_h_r_24_34990 = net_34990;
  assign seg_10_11_sp4_h_r_30_34998 = net_34998;
  assign seg_10_11_sp4_r_v_b_6_42302 = seg_11_9_sp4_v_b_30_42302;
  assign seg_10_11_sp4_v_b_3_38466 = seg_10_10_sp4_v_b_14_38466;
  assign seg_10_12_sp12_v_b_0_41270 = seg_10_4_sp12_v_b_16_41270;
  assign seg_10_12_sp4_h_r_20_38955 = net_38955;
  assign seg_10_12_sp4_v_b_0_38588 = seg_9_11_sp4_r_v_b_13_38588;
  assign seg_10_12_sp4_v_b_7_38593 = seg_9_10_sp4_r_v_b_31_38593;
  assign seg_10_12_sp4_v_b_8_38596 = seg_10_10_sp4_v_b_32_38596;
  assign seg_10_13_lutff_1_out_38933 = net_38933;
  assign seg_10_13_lutff_2_out_38934 = net_38934;
  assign seg_10_14_sp4_h_l_46_28036 = seg_7_14_sp4_h_r_22_28036;
  assign seg_10_14_sp4_h_r_10_43023 = net_43023;
  assign seg_10_14_sp4_h_r_16_39197 = net_39197;
  assign seg_10_14_sp4_h_r_24_35359 = net_35359;
  assign seg_10_14_sp4_r_v_b_19_42794 = net_42794;
  assign seg_10_14_sp4_r_v_b_23_42798 = net_42798;
  assign seg_10_14_sp4_v_b_14_38958 = net_38958;
  assign seg_10_15_lutff_0_out_39178 = net_39178;
  assign seg_10_15_lutff_4_out_39182 = net_39182;
  assign seg_10_15_lutff_7_out_39185 = net_39185;
  assign seg_10_15_neigh_op_bnl_2_35226 = seg_9_14_lutff_2_out_35226;
  assign seg_10_15_sp4_h_l_36_28136 = seg_9_15_sp4_h_r_36_28136;
  assign seg_10_15_sp4_h_r_10_43146 = seg_12_15_sp4_h_r_34_43146;
  assign seg_10_15_sp4_v_b_36_39325 = net_39325;
  assign seg_10_15_sp4_v_b_3_38958 = seg_10_14_sp4_v_b_14_38958;
  assign seg_10_16_lutff_0_out_39301 = net_39301;
  assign seg_10_16_lutff_1_out_39302 = net_39302;
  assign seg_10_16_lutff_3_out_39304 = net_39304;
  assign seg_10_16_lutff_4_out_39305 = net_39305;
  assign seg_10_16_lutff_5_out_39306 = net_39306;
  assign seg_10_16_sp4_h_r_3_43272 = seg_13_16_sp4_h_r_38_43272;
  assign seg_10_16_sp4_h_r_7_43276 = seg_11_16_sp4_h_r_18_43276;
  assign seg_10_16_sp4_v_t_46_39581 = seg_9_18_sp4_r_v_b_35_39581;
  assign seg_10_17_lutff_0_out_39424 = net_39424;
  assign seg_10_17_lutff_1_out_39425 = net_39425;
  assign seg_10_17_lutff_2_out_39426 = net_39426;
  assign seg_10_17_lutff_4_out_39428 = net_39428;
  assign seg_10_17_lutff_6_out_39430 = net_39430;
  assign seg_10_17_lutff_7_out_39431 = net_39431;
  assign seg_10_17_neigh_op_bot_0_39301 = seg_10_16_lutff_0_out_39301;
  assign seg_10_17_neigh_op_bot_4_39305 = seg_10_16_lutff_4_out_39305;
  assign seg_10_17_neigh_op_bot_5_39306 = seg_10_16_lutff_5_out_39306;
  assign seg_10_17_neigh_op_rgt_3_43258 = seg_11_17_lutff_3_out_43258;
  assign seg_10_17_neigh_op_rgt_4_43259 = seg_11_17_lutff_4_out_43259;
  assign seg_10_17_neigh_op_rgt_7_43262 = seg_11_17_lutff_7_out_43262;
  assign seg_10_17_sp4_h_r_11_43393 = seg_13_17_sp4_h_r_46_43393;
  assign seg_10_18_lutff_1_out_39548 = net_39548;
  assign seg_10_18_lutff_2_out_39549 = net_39549;
  assign seg_10_18_lutff_3_out_39550 = net_39550;
  assign seg_10_18_lutff_5_out_39552 = net_39552;
  assign seg_10_18_lutff_6_out_39553 = net_39553;
  assign seg_10_18_lutff_7_out_39554 = net_39554;
  assign seg_10_18_neigh_op_lft_0_35716 = seg_9_18_lutff_0_out_35716;
  assign seg_10_18_neigh_op_lft_2_35718 = seg_9_18_lutff_2_out_35718;
  assign seg_10_18_neigh_op_lft_5_35721 = seg_9_18_lutff_5_out_35721;
  assign seg_10_18_neigh_op_lft_6_35722 = seg_9_18_lutff_6_out_35722;
  assign seg_10_18_neigh_op_lft_7_35723 = seg_9_18_lutff_7_out_35723;
  assign seg_10_18_neigh_op_rgt_1_43379 = seg_11_18_lutff_1_out_43379;
  assign seg_10_18_sp4_h_r_0_43513 = net_43513;
  assign seg_10_18_sp4_h_r_3_43518 = seg_13_18_sp4_h_r_38_43518;
  assign seg_10_18_sp4_h_r_8_43523 = net_43523;
  assign seg_10_18_sp4_r_v_b_8_43165 = seg_11_16_sp4_v_b_32_43165;
  assign seg_10_19_neigh_op_rgt_1_43502 = seg_11_19_lutff_1_out_43502;
  assign seg_10_19_sp12_v_b_2_42281 = seg_10_9_sp12_v_b_22_42281;
  assign seg_10_19_sp4_r_v_b_15_43405 = net_43405;
  assign seg_10_19_sp4_r_v_b_3_43281 = net_43281;
  assign seg_10_1_lutff_1_out_37416 = net_37416;
  assign seg_10_1_lutff_2_out_37417 = net_37417;
  assign seg_10_1_lutff_5_out_37420 = net_37420;
  assign seg_10_1_lutff_6_out_37421 = net_37421;
  assign seg_10_1_lutff_7_out_37422 = net_37422;
  assign seg_10_1_neigh_op_lft_1_33585 = seg_9_1_lutff_1_out_33585;
  assign seg_10_1_neigh_op_lft_3_33587 = seg_9_1_lutff_3_out_33587;
  assign seg_10_1_neigh_op_lft_4_33588 = seg_9_1_lutff_4_out_33588;
  assign seg_10_1_neigh_op_lft_6_33590 = seg_9_1_lutff_6_out_33590;
  assign seg_10_1_neigh_op_top_5_37548 = seg_10_2_lutff_5_out_37548;
  assign seg_10_1_neigh_op_top_7_37550 = seg_10_2_lutff_7_out_37550;
  assign seg_10_1_sp4_h_r_9_41397 = seg_13_1_sp4_h_r_44_41397;
  assign seg_10_1_sp4_r_v_b_47_41440 = net_41440;
  assign seg_10_2_lutff_0_out_37543 = net_37543;
  assign seg_10_2_lutff_1_out_37544 = net_37544;
  assign seg_10_2_lutff_2_out_37545 = net_37545;
  assign seg_10_2_lutff_3_out_37546 = net_37546;
  assign seg_10_2_lutff_4_out_37547 = net_37547;
  assign seg_10_2_lutff_5_out_37548 = net_37548;
  assign seg_10_2_lutff_6_out_37549 = net_37549;
  assign seg_10_2_lutff_7_out_37550 = net_37550;
  assign seg_10_2_sp4_h_r_28_33889 = seg_8_2_sp4_h_r_4_33889;
  assign seg_10_2_sp4_v_b_39_37729 = seg_10_5_sp4_v_b_2_37729;
  assign seg_10_2_sp4_v_t_44_37857 = seg_9_6_sp4_r_v_b_9_37857;
  assign seg_10_3_lutff_0_out_37702 = net_37702;
  assign seg_10_3_lutff_1_out_37703 = net_37703;
  assign seg_10_3_lutff_2_out_37704 = net_37704;
  assign seg_10_3_lutff_3_out_37705 = net_37705;
  assign seg_10_3_lutff_4_out_37706 = net_37706;
  assign seg_10_3_lutff_5_out_37707 = net_37707;
  assign seg_10_3_lutff_6_out_37708 = net_37708;
  assign seg_10_3_lutff_7_out_37709 = net_37709;
  assign seg_10_3_sp4_h_l_46_26914 = seg_7_3_sp4_h_r_22_26914;
  assign seg_10_3_sp4_h_r_0_41668 = seg_12_3_sp4_h_r_24_41668;
  assign seg_10_3_sp4_h_r_37_30175 = seg_7_3_sp4_h_r_0_30175;
  assign seg_10_3_sp4_h_r_45_30185 = seg_7_3_sp4_h_r_8_30185;
  assign seg_10_3_sp4_v_b_12_37597 = net_37597;
  assign seg_10_3_sp4_v_b_36_37849 = seg_10_5_sp4_v_b_12_37849;
  assign seg_10_3_sp4_v_t_47_37983 = seg_10_7_sp4_v_b_10_37983;
  assign seg_10_4_lutff_1_out_37826 = net_37826;
  assign seg_10_4_lutff_3_out_37828 = net_37828;
  assign seg_10_4_lutff_6_out_37831 = net_37831;
  assign seg_10_4_neigh_op_lft_6_34000 = seg_9_4_lutff_6_out_34000;
  assign seg_10_4_neigh_op_lft_7_34001 = seg_9_4_lutff_7_out_34001;
  assign seg_10_4_sp12_v_b_16_41270 = net_41270;
  assign seg_10_4_sp4_h_r_10_41793 = net_41793;
  assign seg_10_4_sp4_h_r_1_41792 = seg_13_4_sp4_h_r_36_41792;
  assign seg_10_4_sp4_h_r_3_41796 = seg_13_4_sp4_h_r_38_41796;
  assign seg_10_4_sp4_r_v_b_31_41686 = net_41686;
  assign seg_10_4_sp4_v_b_1_37597 = seg_10_3_sp4_v_b_12_37597;
  assign seg_10_5_lutff_4_out_37952 = net_37952;
  assign seg_10_5_lutff_5_out_37953 = net_37953;
  assign seg_10_5_lutff_7_out_37955 = net_37955;
  assign seg_10_5_neigh_op_lft_0_34117 = seg_9_5_lutff_0_out_34117;
  assign seg_10_5_neigh_op_tnl_2_34242 = seg_9_6_lutff_2_out_34242;
  assign seg_10_5_sp4_v_b_12_37849 = net_37849;
  assign seg_10_5_sp4_v_b_2_37729 = net_37729;
  assign seg_10_6_neigh_op_bnr_2_41781 = seg_11_5_lutff_2_out_41781;
  assign seg_10_6_neigh_op_rgt_1_41903 = seg_11_6_lutff_1_out_41903;
  assign seg_10_6_sp4_h_r_24_34375 = net_34375;
  assign seg_10_6_sp4_h_r_2_42041 = net_42041;
  assign seg_10_6_sp4_v_b_30_38102 = net_38102;
  assign seg_10_7_lutff_0_out_38194 = net_38194;
  assign seg_10_7_lutff_1_out_38195 = net_38195;
  assign seg_10_7_lutff_3_out_38197 = net_38197;
  assign seg_10_7_lutff_7_out_38201 = net_38201;
  assign seg_10_7_neigh_op_lft_0_34363 = seg_9_7_lutff_0_out_34363;
  assign seg_10_7_neigh_op_tnl_3_34489 = seg_9_8_lutff_3_out_34489;
  assign seg_10_7_neigh_op_top_4_38321 = seg_10_8_lutff_4_out_38321;
  assign seg_10_7_sp12_h_r_0_42156 = seg_18_7_sp12_h_r_16_42156;
  assign seg_10_7_sp4_h_r_16_38336 = net_38336;
  assign seg_10_7_sp4_h_r_24_34498 = net_34498;
  assign seg_10_7_sp4_r_v_b_33_42057 = net_42057;
  assign seg_10_7_sp4_v_b_10_37983 = net_37983;
  assign seg_10_7_sp4_v_b_24_38219 = net_38219;
  assign seg_10_7_sp4_v_b_3_37974 = seg_9_7_sp4_r_v_b_3_37974;
  assign seg_10_7_sp4_v_b_41_38346 = seg_10_10_sp4_v_b_4_38346;
  assign seg_10_7_sp4_v_t_36_38464 = seg_9_11_sp4_r_v_b_1_38464;
  assign seg_10_8_lutff_1_out_38318 = net_38318;
  assign seg_10_8_lutff_3_out_38320 = net_38320;
  assign seg_10_8_lutff_4_out_38321 = net_38321;
  assign seg_10_8_lutff_5_out_38322 = net_38322;
  assign seg_10_8_lutff_6_out_38323 = net_38323;
  assign seg_10_8_lutff_7_out_38324 = net_38324;
  assign seg_10_8_neigh_op_lft_2_34488 = seg_9_8_lutff_2_out_34488;
  assign seg_10_8_neigh_op_lft_4_34490 = seg_9_8_lutff_4_out_34490;
  assign seg_10_8_neigh_op_lft_5_34491 = seg_9_8_lutff_5_out_34491;
  assign seg_10_8_neigh_op_lft_6_34492 = seg_9_8_lutff_6_out_34492;
  assign seg_10_8_neigh_op_tnl_0_34609 = seg_9_9_lutff_0_out_34609;
  assign seg_10_8_sp4_h_r_14_38457 = net_38457;
  assign seg_10_8_sp4_h_r_46_30793 = net_30793;
  assign seg_10_8_sp4_r_v_b_1_41926 = net_41926;
  assign seg_10_8_sp4_r_v_b_47_42306 = net_42306;
  assign seg_10_8_sp4_v_b_6_38102 = seg_10_6_sp4_v_b_30_38102;
  assign seg_10_8_sp4_v_t_37_38588 = seg_9_11_sp4_r_v_b_13_38588;
  assign seg_10_8_sp4_v_t_41_38592 = seg_9_11_sp4_r_v_b_17_38592;
  assign seg_10_9_neigh_op_bot_7_38324 = seg_10_8_lutff_7_out_38324;
  assign seg_10_9_sp12_v_b_22_42281 = net_42281;
  assign seg_10_9_sp4_v_b_0_38219 = seg_10_7_sp4_v_b_24_38219;
  assign seg_10_9_sp4_v_b_11_38228 = seg_9_7_sp4_r_v_b_35_38228;
  assign seg_11_10_lutff_1_out_42395 = net_42395;
  assign seg_11_10_lutff_4_out_42398 = net_42398;
  assign seg_11_10_lutff_7_out_42401 = net_42401;
  assign seg_11_10_neigh_op_bot_7_42278 = seg_11_9_lutff_7_out_42278;
  assign seg_11_10_neigh_op_rgt_1_46226 = seg_12_10_lutff_1_out_46226;
  assign seg_11_10_sp4_h_r_3_46365 = seg_12_10_sp4_h_r_14_46365;
  assign seg_11_10_sp4_h_r_7_46369 = seg_12_10_sp4_h_r_18_46369;
  assign seg_11_11_lutff_1_out_42518 = net_42518;
  assign seg_11_11_lutff_4_out_42521 = net_42521;
  assign seg_11_11_lutff_5_out_42522 = net_42522;
  assign seg_11_11_lutff_6_out_42523 = net_42523;
  assign seg_11_11_neigh_op_bot_4_42398 = seg_11_10_lutff_4_out_42398;
  assign seg_11_11_neigh_op_lft_6_38692 = seg_10_11_lutff_6_out_38692;
  assign seg_11_11_sp12_h_r_22_2407 = net_2407;
  assign seg_11_11_sp12_v_b_22_46358 = net_46358;
  assign seg_11_11_sp12_v_b_4_45216 = net_45216;
  assign seg_11_11_sp4_h_l_38_31164 = seg_8_11_sp4_h_r_14_31164;
  assign seg_11_11_sp4_h_l_41_31165 = seg_9_11_sp4_h_r_28_31165;
  assign seg_11_11_sp4_h_r_16_42659 = net_42659;
  assign seg_11_11_sp4_r_v_b_15_46252 = net_46252;
  assign seg_11_11_sp4_r_v_b_21_46258 = net_46258;
  assign seg_11_11_sp4_r_v_b_23_46260 = net_46260;
  assign seg_11_11_sp4_r_v_b_44_46503 = seg_12_13_sp4_v_b_20_46503;
  assign seg_11_11_sp4_v_b_0_42296 = seg_11_9_sp4_v_b_24_42296;
  assign seg_11_11_sp4_v_b_10_42306 = seg_10_8_sp4_r_v_b_47_42306;
  assign seg_11_11_sp4_v_b_6_42302 = seg_11_9_sp4_v_b_30_42302;
  assign seg_11_12_lutff_2_out_42642 = net_42642;
  assign seg_11_12_neigh_op_bnl_1_38687 = seg_10_11_lutff_1_out_38687;
  assign seg_11_12_neigh_op_rgt_0_46471 = seg_12_12_lutff_0_out_46471;
  assign seg_11_12_neigh_op_tnr_2_46596 = seg_12_13_lutff_2_out_46596;
  assign seg_11_12_sp12_v_b_10_45743 = net_45743;
  assign seg_11_12_sp4_h_r_10_46608 = seg_13_12_sp4_h_r_34_46608;
  assign seg_11_12_sp4_h_r_2_46610 = net_46610;
  assign seg_11_12_sp4_r_v_b_1_46249 = net_46249;
  assign seg_11_12_sp4_r_v_b_24_46496 = seg_12_14_sp4_v_b_0_46496;
  assign seg_11_12_sp4_v_b_40_42791 = net_42791;
  assign seg_11_13_lutff_4_out_42767 = net_42767;
  assign seg_11_13_sp12_v_b_0_45216 = seg_11_11_sp12_v_b_4_45216;
  assign seg_11_13_sp12_v_b_1_45215 = seg_11_8_sp12_v_b_10_45215;
  assign seg_11_13_sp4_h_r_11_46732 = seg_14_13_sp4_h_r_46_46732;
  assign seg_11_13_sp4_h_r_1_46730 = seg_14_13_sp4_h_r_36_46730;
  assign seg_11_13_sp4_h_r_25_39068 = seg_12_13_sp4_h_r_36_39068;
  assign seg_11_13_sp4_h_r_34_39069 = seg_9_13_sp4_h_r_10_39069;
  assign seg_11_13_sp4_h_r_9_46740 = seg_12_13_sp4_h_r_20_46740;
  assign seg_11_13_sp4_v_b_20_42672 = net_42672;
  assign seg_11_14_neigh_op_tnr_3_46843 = seg_12_15_lutff_3_out_46843;
  assign seg_11_14_sp12_v_b_14_46235 = net_46235;
  assign seg_11_14_sp12_v_b_8_45867 = net_45867;
  assign seg_11_14_sp4_h_l_39_31532 = seg_9_14_sp4_h_r_26_31532;
  assign seg_11_14_sp4_h_r_0_46852 = net_46852;
  assign seg_11_14_sp4_h_r_10_46854 = seg_13_14_sp4_h_r_34_46854;
  assign seg_11_14_sp4_h_r_42_35368 = net_35368;
  assign seg_11_14_sp4_h_r_4_46858 = seg_13_14_sp4_h_r_28_46858;
  assign seg_11_14_sp4_r_v_b_21_46627 = net_46627;
  assign seg_11_14_sp4_v_b_9_42672 = seg_11_13_sp4_v_b_20_42672;
  assign seg_11_15_lutff_0_out_43009 = net_43009;
  assign seg_11_15_lutff_6_out_43015 = net_43015;
  assign seg_11_15_neigh_op_rgt_2_46842 = seg_12_15_lutff_2_out_46842;
  assign seg_11_15_sp4_h_l_36_31652 = seg_8_15_sp4_h_r_12_31652;
  assign seg_11_15_sp4_h_r_46_35485 = net_35485;
  assign seg_11_15_sp4_h_r_9_46986 = seg_12_15_sp4_h_r_20_46986;
  assign seg_11_15_sp4_r_v_b_12_46741 = seg_12_13_sp4_v_b_36_46741;
  assign seg_11_15_sp4_v_b_10_42798 = seg_10_14_sp4_r_v_b_23_42798;
  assign seg_11_15_sp4_v_b_24_43034 = net_43034;
  assign seg_11_15_sp4_v_b_34_43044 = net_43044;
  assign seg_11_15_sp4_v_b_36_43156 = net_43156;
  assign seg_11_15_sp4_v_b_5_42791 = seg_11_12_sp4_v_b_40_42791;
  assign seg_11_15_sp4_v_b_6_42794 = seg_10_14_sp4_r_v_b_19_42794;
  assign seg_11_15_sp4_v_t_38_43281 = seg_10_19_sp4_r_v_b_3_43281;
  assign seg_11_16_lutff_3_out_43135 = net_43135;
  assign seg_11_16_lutff_4_out_43136 = net_43136;
  assign seg_11_16_sp12_v_b_2_45743 = seg_11_12_sp12_v_b_10_45743;
  assign seg_11_16_sp4_h_r_18_43276 = net_43276;
  assign seg_11_16_sp4_r_v_b_45_47119 = seg_11_18_sp4_r_v_b_21_47119;
  assign seg_11_16_sp4_v_b_32_43165 = net_43165;
  assign seg_11_16_sp4_v_t_39_43405 = seg_10_19_sp4_r_v_b_15_43405;
  assign seg_11_17_lutff_0_out_43255 = net_43255;
  assign seg_11_17_lutff_2_out_43257 = net_43257;
  assign seg_11_17_lutff_3_out_43258 = net_43258;
  assign seg_11_17_lutff_4_out_43259 = net_43259;
  assign seg_11_17_lutff_5_out_43260 = net_43260;
  assign seg_11_17_lutff_6_out_43261 = net_43261;
  assign seg_11_17_lutff_7_out_43262 = net_43262;
  assign seg_11_17_sp4_h_r_22_43393 = seg_13_17_sp4_h_r_46_43393;
  assign seg_11_17_sp4_h_r_6_47229 = seg_13_17_sp4_h_r_30_47229;
  assign seg_11_17_sp4_r_v_b_10_46875 = seg_12_15_sp4_v_b_34_46875;
  assign seg_11_17_sp4_v_b_0_43034 = seg_11_15_sp4_v_b_24_43034;
  assign seg_11_17_sp4_v_b_10_43044 = seg_11_15_sp4_v_b_34_43044;
  assign seg_11_18_lutff_1_out_43379 = net_43379;
  assign seg_11_18_neigh_op_bot_5_43260 = seg_11_17_lutff_5_out_43260;
  assign seg_11_18_neigh_op_bot_6_43261 = seg_11_17_lutff_6_out_43261;
  assign seg_11_18_neigh_op_rgt_2_47211 = seg_12_18_lutff_2_out_47211;
  assign seg_11_18_neigh_op_rgt_4_47213 = seg_12_18_lutff_4_out_47213;
  assign seg_11_18_neigh_op_tnr_3_47335 = seg_12_19_lutff_3_out_47335;
  assign seg_11_18_sp12_v_b_0_45867 = seg_11_14_sp12_v_b_8_45867;
  assign seg_11_18_sp12_v_b_6_46235 = seg_11_14_sp12_v_b_14_46235;
  assign seg_11_18_sp4_r_v_b_15_47113 = net_47113;
  assign seg_11_18_sp4_r_v_b_21_47119 = net_47119;
  assign seg_11_18_sp4_r_v_b_27_47235 = net_47235;
  assign seg_11_18_sp4_v_b_1_43156 = seg_11_15_sp4_v_b_36_43156;
  assign seg_11_19_lutff_1_out_43502 = net_43502;
  assign seg_11_1_sp4_r_v_b_9_45276 = net_45276;
  assign seg_11_22_sp12_v_b_1_46358 = seg_11_11_sp12_v_b_22_46358;
  assign seg_11_2_lutff_2_out_41376 = net_41376;
  assign seg_11_2_lutff_4_out_41378 = net_41378;
  assign seg_11_2_lutff_7_out_41381 = net_41381;
  assign seg_11_2_neigh_op_bnl_1_37416 = seg_10_1_lutff_1_out_37416;
  assign seg_11_2_neigh_op_bnl_2_37417 = seg_10_1_lutff_2_out_37417;
  assign seg_11_2_neigh_op_bnl_7_37422 = seg_10_1_lutff_7_out_37422;
  assign seg_11_2_neigh_op_bnr_1_45078 = seg_12_1_lutff_1_out_45078;
  assign seg_11_2_neigh_op_rgt_3_45208 = seg_12_2_lutff_3_out_45208;
  assign seg_11_2_sp4_h_r_10_45378 = net_45378;
  assign seg_11_2_sp4_h_r_28_37720 = net_37720;
  assign seg_11_2_sp4_h_r_34_37716 = net_37716;
  assign seg_11_2_sp4_v_b_26_41431 = seg_11_4_sp4_v_b_2_41431;
  assign seg_11_2_sp4_v_b_37_41558 = seg_11_5_sp4_v_b_0_41558;
  assign seg_11_2_sp4_v_b_38_41559 = seg_11_4_sp4_v_b_14_41559;
  assign seg_11_2_sp4_v_b_39_41560 = seg_11_5_sp4_v_b_2_41560;
  assign seg_11_3_lutff_1_out_41534 = net_41534;
  assign seg_11_3_lutff_2_out_41535 = net_41535;
  assign seg_11_3_lutff_3_out_41536 = net_41536;
  assign seg_11_3_lutff_4_out_41537 = net_41537;
  assign seg_11_3_lutff_5_out_41538 = net_41538;
  assign seg_11_3_lutff_6_out_41539 = net_41539;
  assign seg_11_3_lutff_7_out_41540 = net_41540;
  assign seg_11_3_neigh_op_bnl_1_37544 = seg_10_2_lutff_1_out_37544;
  assign seg_11_3_neigh_op_bnl_4_37547 = seg_10_2_lutff_4_out_37547;
  assign seg_11_3_neigh_op_bot_7_41381 = seg_11_2_lutff_7_out_41381;
  assign seg_11_3_neigh_op_lft_0_37702 = seg_10_3_lutff_0_out_37702;
  assign seg_11_3_neigh_op_lft_1_37703 = seg_10_3_lutff_1_out_37703;
  assign seg_11_3_neigh_op_lft_2_37704 = seg_10_3_lutff_2_out_37704;
  assign seg_11_3_neigh_op_lft_3_37705 = seg_10_3_lutff_3_out_37705;
  assign seg_11_3_neigh_op_lft_4_37706 = seg_10_3_lutff_4_out_37706;
  assign seg_11_3_neigh_op_lft_5_37707 = seg_10_3_lutff_5_out_37707;
  assign seg_11_3_neigh_op_lft_6_37708 = seg_10_3_lutff_6_out_37708;
  assign seg_11_3_neigh_op_lft_7_37709 = seg_10_3_lutff_7_out_37709;
  assign seg_11_3_sp4_v_b_30_41564 = seg_11_5_sp4_v_b_6_41564;
  assign seg_11_3_sp4_v_b_32_41566 = seg_11_5_sp4_v_b_8_41566;
  assign seg_11_3_sp4_v_b_38_41682 = seg_11_5_sp4_v_b_14_41682;
  assign seg_11_4_lutff_3_out_41659 = net_41659;
  assign seg_11_4_lutff_5_out_41661 = net_41661;
  assign seg_11_4_neigh_op_bot_1_41534 = seg_11_3_lutff_1_out_41534;
  assign seg_11_4_neigh_op_bot_2_41535 = seg_11_3_lutff_2_out_41535;
  assign seg_11_4_neigh_op_bot_3_41536 = seg_11_3_lutff_3_out_41536;
  assign seg_11_4_neigh_op_bot_4_41537 = seg_11_3_lutff_4_out_41537;
  assign seg_11_4_neigh_op_bot_5_41538 = seg_11_3_lutff_5_out_41538;
  assign seg_11_4_neigh_op_bot_6_41539 = seg_11_3_lutff_6_out_41539;
  assign seg_11_4_neigh_op_bot_7_41540 = seg_11_3_lutff_7_out_41540;
  assign seg_11_4_neigh_op_rgt_5_45492 = seg_12_4_lutff_5_out_45492;
  assign seg_11_4_sp12_h_r_6_34126 = net_34126;
  assign seg_11_4_sp4_h_l_40_30305 = seg_8_4_sp4_h_r_16_30305;
  assign seg_11_4_sp4_h_l_46_30301 = seg_8_4_sp4_h_r_22_30301;
  assign seg_11_4_sp4_h_r_1_45623 = seg_14_4_sp4_h_r_36_45623;
  assign seg_11_4_sp4_h_r_28_37966 = net_37966;
  assign seg_11_4_sp4_h_r_3_45627 = seg_12_4_sp4_h_r_14_45627;
  assign seg_11_4_sp4_h_r_7_45631 = seg_12_4_sp4_h_r_18_45631;
  assign seg_11_4_sp4_h_r_8_45632 = net_45632;
  assign seg_11_4_sp4_r_v_b_5_45264 = net_45264;
  assign seg_11_4_sp4_v_b_10_41440 = seg_10_1_sp4_r_v_b_47_41440;
  assign seg_11_4_sp4_v_b_14_41559 = net_41559;
  assign seg_11_4_sp4_v_b_2_41431 = net_41431;
  assign seg_11_4_sp4_v_t_36_41926 = seg_10_8_sp4_r_v_b_1_41926;
  assign seg_11_4_sp4_v_t_41_41931 = seg_11_8_sp4_v_b_4_41931;
  assign seg_11_5_lutff_2_out_41781 = net_41781;
  assign seg_11_5_lutff_3_out_41782 = net_41782;
  assign seg_11_5_lutff_6_out_41785 = net_41785;
  assign seg_11_5_neigh_op_bot_3_41659 = seg_11_4_lutff_3_out_41659;
  assign seg_11_5_neigh_op_lft_7_37955 = seg_10_5_lutff_7_out_37955;
  assign seg_11_5_neigh_op_top_4_41906 = seg_11_6_lutff_4_out_41906;
  assign seg_11_5_neigh_op_top_7_41909 = seg_11_6_lutff_7_out_41909;
  assign seg_11_5_sp4_h_r_10_45747 = net_45747;
  assign seg_11_5_sp4_h_r_26_38087 = net_38087;
  assign seg_11_5_sp4_h_r_4_45751 = net_45751;
  assign seg_11_5_sp4_r_v_b_43_45764 = net_45764;
  assign seg_11_5_sp4_v_b_0_41558 = net_41558;
  assign seg_11_5_sp4_v_b_14_41682 = net_41682;
  assign seg_11_5_sp4_v_b_20_41688 = net_41688;
  assign seg_11_5_sp4_v_b_2_41560 = net_41560;
  assign seg_11_5_sp4_v_b_6_41564 = net_41564;
  assign seg_11_5_sp4_v_b_8_41566 = net_41566;
  assign seg_11_5_sp4_v_t_44_42057 = seg_10_7_sp4_r_v_b_33_42057;
  assign seg_11_6_lutff_0_out_41902 = net_41902;
  assign seg_11_6_lutff_1_out_41903 = net_41903;
  assign seg_11_6_lutff_4_out_41906 = net_41906;
  assign seg_11_6_lutff_7_out_41909 = net_41909;
  assign seg_11_6_neigh_op_tnl_1_38195 = seg_10_7_lutff_1_out_38195;
  assign seg_11_6_neigh_op_tnl_3_38197 = seg_10_7_lutff_3_out_38197;
  assign seg_11_6_sp4_h_r_18_42046 = net_42046;
  assign seg_11_6_sp4_h_r_2_45872 = net_45872;
  assign seg_11_6_sp4_h_r_46_34378 = seg_9_6_sp4_h_r_22_34378;
  assign seg_11_6_sp4_r_v_b_35_45767 = net_45767;
  assign seg_11_6_sp4_v_b_7_41686 = seg_10_4_sp4_r_v_b_31_41686;
  assign seg_11_6_sp4_v_b_9_41688 = seg_11_5_sp4_v_b_20_41688;
  assign seg_11_7_neigh_op_lft_0_38194 = seg_10_7_lutff_0_out_38194;
  assign seg_11_7_sp12_h_r_1_45988 = seg_18_7_sp12_h_r_14_45988;
  assign seg_11_7_sp4_h_r_0_45991 = net_45991;
  assign seg_11_7_sp4_h_r_10_45993 = net_45993;
  assign seg_11_7_sp4_h_r_11_45994 = seg_12_7_sp4_h_r_22_45994;
  assign seg_11_7_sp4_h_r_3_45996 = seg_14_7_sp4_h_r_38_45996;
  assign seg_11_7_sp4_r_v_b_41_46008 = net_46008;
  assign seg_11_8_lutff_0_out_42148 = net_42148;
  assign seg_11_8_lutff_1_out_42149 = net_42149;
  assign seg_11_8_lutff_2_out_42150 = net_42150;
  assign seg_11_8_lutff_4_out_42152 = net_42152;
  assign seg_11_8_neigh_op_lft_3_38320 = seg_10_8_lutff_3_out_38320;
  assign seg_11_8_neigh_op_lft_6_38323 = seg_10_8_lutff_6_out_38323;
  assign seg_11_8_sp12_h_r_14_19925 = net_19925;
  assign seg_11_8_sp12_h_r_20_7898 = net_7898;
  assign seg_11_8_sp12_h_r_22_1764 = net_1764;
  assign seg_11_8_sp12_v_b_10_45215 = net_45215;
  assign seg_11_8_sp4_h_l_43_30798 = seg_9_8_sp4_h_r_30_30798;
  assign seg_11_8_sp4_h_l_46_30793 = seg_10_8_sp4_h_r_46_30793;
  assign seg_11_8_sp4_h_r_0_46114 = seg_13_8_sp4_h_r_24_46114;
  assign seg_11_8_sp4_h_r_11_46117 = seg_14_8_sp4_h_r_46_46117;
  assign seg_11_8_sp4_h_r_20_42294 = net_42294;
  assign seg_11_8_sp4_h_r_38_34626 = net_34626;
  assign seg_11_8_sp4_h_r_3_46119 = seg_14_8_sp4_h_r_38_46119;
  assign seg_11_8_sp4_h_r_42_34630 = net_34630;
  assign seg_11_8_sp4_h_r_44_34632 = net_34632;
  assign seg_11_8_sp4_h_r_46_34624 = net_34624;
  assign seg_11_8_sp4_h_r_5_46121 = seg_14_8_sp4_h_r_40_46121;
  assign seg_11_8_sp4_r_v_b_17_45885 = net_45885;
  assign seg_11_8_sp4_r_v_b_21_45889 = net_45889;
  assign seg_11_8_sp4_r_v_b_33_46011 = net_46011;
  assign seg_11_8_sp4_v_b_4_41931 = net_41931;
  assign seg_11_9_lutff_1_out_42272 = net_42272;
  assign seg_11_9_lutff_7_out_42278 = net_42278;
  assign seg_11_9_sp12_h_r_3_42402 = seg_16_9_sp12_h_r_12_42402;
  assign seg_11_9_sp4_v_b_24_42296 = net_42296;
  assign seg_11_9_sp4_v_b_30_42302 = net_42302;
  assign seg_12_0_logic_op_tnr_5_48913 = seg_13_1_lutff_5_out_48913;
  assign seg_12_10_lutff_1_out_46226 = net_46226;
  assign seg_12_10_sp12_v_b_1_48926 = seg_12_3_sp12_v_b_14_48926;
  assign seg_12_10_sp4_h_r_14_46365 = net_46365;
  assign seg_12_10_sp4_h_r_18_46369 = net_46369;
  assign seg_12_10_sp4_h_r_46_38701 = net_38701;
  assign seg_12_10_sp4_r_v_b_31_50086 = net_50086;
  assign seg_12_10_sp4_r_v_b_39_50206 = net_50206;
  assign seg_12_10_sp4_r_v_b_45_50212 = net_50212;
  assign seg_12_10_sp4_r_v_b_47_50214 = net_50214;
  assign seg_12_10_sp4_v_b_18_46132 = net_46132;
  assign seg_12_10_sp4_v_b_24_46250 = net_46250;
  assign seg_12_10_sp4_v_b_40_46376 = net_46376;
  assign seg_12_10_sp4_v_b_8_46012 = net_46012;
  assign seg_12_11_sp4_h_l_36_34991 = seg_9_11_sp4_h_r_12_34991;
  assign seg_12_11_sp4_h_r_4_50320 = net_50320;
  assign seg_12_11_sp4_h_r_7_50323 = seg_15_11_sp4_h_r_42_50323;
  assign seg_12_11_sp4_r_v_b_23_50091 = net_50091;
  assign seg_12_11_sp4_r_v_b_41_50331 = net_50331;
  assign seg_12_11_sp4_r_v_b_43_50333 = net_50333;
  assign seg_12_11_sp4_r_v_b_45_50335 = net_50335;
  assign seg_12_11_sp4_v_b_11_46136 = seg_12_8_sp4_v_b_46_46136;
  assign seg_12_11_sp4_v_b_7_46132 = seg_12_10_sp4_v_b_18_46132;
  assign seg_12_11_sp4_v_t_39_46621 = seg_12_15_sp4_v_b_2_46621;
  assign seg_12_12_lutff_0_out_46471 = net_46471;
  assign seg_12_12_lutff_1_out_46472 = net_46472;
  assign seg_12_12_neigh_op_rgt_5_50307 = seg_13_12_lutff_5_out_50307;
  assign seg_12_12_neigh_op_top_2_46596 = seg_12_13_lutff_2_out_46596;
  assign seg_12_12_sp12_v_b_0_48932 = seg_12_6_sp12_v_b_12_48932;
  assign seg_12_12_sp4_h_r_6_50445 = net_50445;
  assign seg_12_12_sp4_v_b_0_46250 = seg_12_10_sp4_v_b_24_46250;
  assign seg_12_12_sp4_v_b_10_46260 = seg_11_11_sp4_r_v_b_23_46260;
  assign seg_12_12_sp4_v_b_2_46252 = seg_11_11_sp4_r_v_b_15_46252;
  assign seg_12_12_sp4_v_b_8_46258 = seg_11_11_sp4_r_v_b_21_46258;
  assign seg_12_12_sp4_v_t_38_46743 = seg_12_15_sp4_v_b_14_46743;
  assign seg_12_12_sp4_v_t_42_46747 = seg_12_15_sp4_v_b_18_46747;
  assign seg_12_12_sp4_v_t_44_46749 = seg_12_15_sp4_v_b_20_46749;
  assign seg_12_13_lutff_0_out_46594 = net_46594;
  assign seg_12_13_lutff_2_out_46596 = net_46596;
  assign seg_12_13_lutff_3_out_46597 = net_46597;
  assign seg_12_13_lutff_4_out_46598 = net_46598;
  assign seg_12_13_lutff_6_out_46600 = net_46600;
  assign seg_12_13_sp4_h_r_20_46740 = net_46740;
  assign seg_12_13_sp4_h_r_36_39068 = net_39068;
  assign seg_12_13_sp4_r_v_b_37_50573 = net_50573;
  assign seg_12_13_sp4_r_v_b_42_50578 = seg_13_15_sp4_v_b_18_50578;
  assign seg_12_13_sp4_r_v_b_43_50579 = net_50579;
  assign seg_12_13_sp4_r_v_b_5_50207 = net_50207;
  assign seg_12_13_sp4_v_b_20_46503 = net_46503;
  assign seg_12_13_sp4_v_b_36_46741 = net_46741;
  assign seg_12_13_sp4_v_b_5_46376 = seg_12_10_sp4_v_b_40_46376;
  assign seg_12_14_lutff_1_out_46718 = net_46718;
  assign seg_12_14_lutff_3_out_46720 = net_46720;
  assign seg_12_14_lutff_4_out_46721 = net_46721;
  assign seg_12_14_lutff_5_out_46722 = net_46722;
  assign seg_12_14_neigh_op_rgt_1_50549 = seg_13_14_lutff_1_out_50549;
  assign seg_12_14_sp4_h_l_37_35359 = seg_10_14_sp4_h_r_24_35359;
  assign seg_12_14_sp4_r_v_b_13_50450 = net_50450;
  assign seg_12_14_sp4_v_b_0_46496 = net_46496;
  assign seg_12_14_sp4_v_b_9_46503 = seg_12_13_sp4_v_b_20_46503;
  assign seg_12_14_sp4_v_t_46_46997 = seg_12_15_sp4_v_b_46_46997;
  assign seg_12_15_lutff_0_out_46840 = net_46840;
  assign seg_12_15_lutff_2_out_46842 = net_46842;
  assign seg_12_15_lutff_3_out_46843 = net_46843;
  assign seg_12_15_lutff_4_out_46844 = net_46844;
  assign seg_12_15_lutff_5_out_46845 = net_46845;
  assign seg_12_15_neigh_op_bnr_2_50550 = seg_13_14_lutff_2_out_50550;
  assign seg_12_15_neigh_op_tnr_3_50797 = seg_13_16_lutff_3_out_50797;
  assign seg_12_15_neigh_op_top_3_46966 = seg_12_16_lutff_3_out_46966;
  assign seg_12_15_sp4_h_l_37_35482 = seg_8_15_sp4_h_r_0_35482;
  assign seg_12_15_sp4_h_l_41_35488 = seg_8_15_sp4_h_r_4_35488;
  assign seg_12_15_sp4_h_r_0_50806 = net_50806;
  assign seg_12_15_sp4_h_r_12_46976 = seg_14_15_sp4_h_r_36_46976;
  assign seg_12_15_sp4_h_r_20_46986 = net_46986;
  assign seg_12_15_sp4_h_r_22_46978 = net_46978;
  assign seg_12_15_sp4_h_r_30_43152 = net_43152;
  assign seg_12_15_sp4_h_r_34_43146 = net_43146;
  assign seg_12_15_sp4_h_r_36_39314 = net_39314;
  assign seg_12_15_sp4_h_r_38_39318 = net_39318;
  assign seg_12_15_sp4_h_r_4_50812 = net_50812;
  assign seg_12_15_sp4_r_v_b_15_50575 = net_50575;
  assign seg_12_15_sp4_r_v_b_19_50579 = seg_12_13_sp4_r_v_b_43_50579;
  assign seg_12_15_sp4_r_v_b_21_50581 = net_50581;
  assign seg_12_15_sp4_r_v_b_23_50583 = net_50583;
  assign seg_12_15_sp4_r_v_b_31_50701 = net_50701;
  assign seg_12_15_sp4_r_v_b_3_50451 = net_50451;
  assign seg_12_15_sp4_r_v_b_5_50453 = net_50453;
  assign seg_12_15_sp4_r_v_b_7_50455 = net_50455;
  assign seg_12_15_sp4_v_b_14_46743 = net_46743;
  assign seg_12_15_sp4_v_b_18_46747 = net_46747;
  assign seg_12_15_sp4_v_b_20_46749 = net_46749;
  assign seg_12_15_sp4_v_b_2_46621 = net_46621;
  assign seg_12_15_sp4_v_b_34_46875 = net_46875;
  assign seg_12_15_sp4_v_b_36_46987 = seg_12_17_sp4_v_b_12_46987;
  assign seg_12_15_sp4_v_b_38_46989 = seg_12_17_sp4_v_b_14_46989;
  assign seg_12_15_sp4_v_b_46_46997 = net_46997;
  assign seg_12_15_sp4_v_b_8_46627 = seg_11_14_sp4_r_v_b_21_46627;
  assign seg_12_15_sp4_v_t_39_47113 = seg_11_18_sp4_r_v_b_15_47113;
  assign seg_12_16_lutff_0_out_46963 = net_46963;
  assign seg_12_16_lutff_1_out_46964 = net_46964;
  assign seg_12_16_lutff_3_out_46966 = net_46966;
  assign seg_12_16_lutff_4_out_46967 = net_46967;
  assign seg_12_16_lutff_5_out_46968 = net_46968;
  assign seg_12_16_lutff_6_out_46969 = net_46969;
  assign seg_12_16_lutff_7_out_46970 = net_46970;
  assign seg_12_16_neigh_op_bot_5_46845 = seg_12_15_lutff_5_out_46845;
  assign seg_12_16_neigh_op_rgt_7_50801 = seg_13_16_lutff_7_out_50801;
  assign seg_12_16_neigh_op_tnr_5_50922 = seg_13_17_lutff_5_out_50922;
  assign seg_12_16_neigh_op_tnr_7_50924 = seg_13_17_lutff_7_out_50924;
  assign seg_12_16_neigh_op_top_1_47087 = seg_12_17_lutff_1_out_47087;
  assign seg_12_16_neigh_op_top_2_47088 = seg_12_17_lutff_2_out_47088;
  assign seg_12_16_neigh_op_top_3_47089 = seg_12_17_lutff_3_out_47089;
  assign seg_12_16_neigh_op_top_6_47092 = seg_12_17_lutff_6_out_47092;
  assign seg_12_16_neigh_op_top_7_47093 = seg_12_17_lutff_7_out_47093;
  assign seg_12_16_sp12_v_b_4_49698 = net_49698;
  assign seg_12_16_sp4_h_r_11_50932 = seg_13_16_sp4_h_r_22_50932;
  assign seg_12_16_sp4_r_v_b_6_50579 = seg_12_13_sp4_r_v_b_43_50579;
  assign seg_12_16_sp4_v_b_1_46741 = seg_12_13_sp4_v_b_36_46741;
  assign seg_12_16_sp4_v_b_9_46749 = seg_12_15_sp4_v_b_20_46749;
  assign seg_12_16_sp4_v_t_38_47235 = seg_11_18_sp4_r_v_b_27_47235;
  assign seg_12_17_lutff_1_out_47087 = net_47087;
  assign seg_12_17_lutff_2_out_47088 = net_47088;
  assign seg_12_17_lutff_3_out_47089 = net_47089;
  assign seg_12_17_lutff_4_out_47090 = net_47090;
  assign seg_12_17_lutff_6_out_47092 = net_47092;
  assign seg_12_17_lutff_7_out_47093 = net_47093;
  assign seg_12_17_neigh_op_bot_0_46963 = seg_12_16_lutff_0_out_46963;
  assign seg_12_17_neigh_op_bot_1_46964 = seg_12_16_lutff_1_out_46964;
  assign seg_12_17_neigh_op_bot_5_46968 = seg_12_16_lutff_5_out_46968;
  assign seg_12_17_sp4_r_v_b_15_50821 = net_50821;
  assign seg_12_17_sp4_v_b_12_46987 = net_46987;
  assign seg_12_17_sp4_v_b_14_46989 = net_46989;
  assign seg_12_18_lutff_2_out_47211 = net_47211;
  assign seg_12_18_lutff_4_out_47213 = net_47213;
  assign seg_12_18_sp4_h_r_3_51180 = seg_13_18_sp4_h_r_14_51180;
  assign seg_12_18_sp4_v_b_11_46997 = seg_12_15_sp4_v_b_46_46997;
  assign seg_12_19_lutff_3_out_47335 = net_47335;
  assign seg_12_1_lutff_1_out_45078 = net_45078;
  assign seg_12_1_lutff_2_out_45079 = net_45079;
  assign seg_12_1_lutff_3_out_45080 = net_45080;
  assign seg_12_1_lutff_4_out_45081 = net_45081;
  assign seg_12_1_neigh_op_tnr_1_49037 = seg_13_2_lutff_1_out_49037;
  assign seg_12_1_sp4_h_r_11_49051 = seg_13_1_sp4_h_r_22_49051;
  assign seg_12_1_sp4_r_v_b_19_49071 = net_49071;
  assign seg_12_1_sp4_r_v_b_21_49074 = net_49074;
  assign seg_12_1_sp4_r_v_b_23_49076 = net_49076;
  assign seg_12_1_sp4_r_v_b_25_49078 = net_49078;
  assign seg_12_1_sp4_r_v_b_35_49089 = net_49089;
  assign seg_12_1_sp4_r_v_b_37_49091 = net_49091;
  assign seg_12_1_sp4_r_v_b_39_49093 = net_49093;
  assign seg_12_1_sp4_r_v_b_41_49096 = net_49096;
  assign seg_12_1_sp4_v_b_34_45257 = net_45257;
  assign seg_12_1_sp4_v_b_9_45276 = seg_11_1_sp4_r_v_b_9_45276;
  assign seg_12_2_lutff_0_out_45205 = net_45205;
  assign seg_12_2_lutff_2_out_45207 = net_45207;
  assign seg_12_2_lutff_3_out_45208 = net_45208;
  assign seg_12_2_lutff_6_out_45211 = net_45211;
  assign seg_12_2_neigh_op_bot_2_45079 = seg_12_1_lutff_2_out_45079;
  assign seg_12_2_neigh_op_bot_3_45080 = seg_12_1_lutff_3_out_45080;
  assign seg_12_2_neigh_op_lft_2_41376 = seg_11_2_lutff_2_out_41376;
  assign seg_12_2_neigh_op_tnr_2_49197 = seg_13_3_lutff_2_out_49197;
  assign seg_12_2_sp4_h_r_2_49211 = net_49211;
  assign seg_12_2_sp4_h_r_38_37719 = net_37719;
  assign seg_12_2_sp4_r_v_b_25_49090 = net_49090;
  assign seg_12_2_sp4_r_v_b_41_49224 = net_49224;
  assign seg_12_2_sp4_v_b_22_45258 = net_45258;
  assign seg_12_2_sp4_v_b_29_45264 = seg_11_4_sp4_r_v_b_5_45264;
  assign seg_12_2_sp4_v_b_34_45271 = net_45271;
  assign seg_12_2_sp4_v_b_38_45390 = net_45390;
  assign seg_12_2_sp4_v_b_40_45392 = net_45392;
  assign seg_12_31_span4_horz_r_6_48880 = net_48880;
  assign seg_12_3_lutff_4_out_45368 = net_45368;
  assign seg_12_3_lutff_5_out_45369 = net_45369;
  assign seg_12_3_lutff_6_out_45370 = net_45370;
  assign seg_12_3_neigh_op_bnl_4_41378 = seg_11_2_lutff_4_out_41378;
  assign seg_12_3_neigh_op_bot_0_45205 = seg_12_2_lutff_0_out_45205;
  assign seg_12_3_neigh_op_bot_2_45207 = seg_12_2_lutff_2_out_45207;
  assign seg_12_3_neigh_op_rgt_6_49201 = seg_13_3_lutff_6_out_49201;
  assign seg_12_3_neigh_op_tnl_5_41661 = seg_11_4_lutff_5_out_41661;
  assign seg_12_3_neigh_op_tnr_6_49324 = seg_13_4_lutff_6_out_49324;
  assign seg_12_3_neigh_op_top_3_45490 = seg_12_4_lutff_3_out_45490;
  assign seg_12_3_sp12_v_b_14_48926 = net_48926;
  assign seg_12_3_sp4_h_r_24_41668 = net_41668;
  assign seg_12_3_sp4_h_r_28_41674 = net_41674;
  assign seg_12_3_sp4_h_r_40_37844 = net_37844;
  assign seg_12_3_sp4_h_r_8_49340 = net_49340;
  assign seg_12_3_sp4_r_v_b_25_49219 = net_49219;
  assign seg_12_3_sp4_r_v_b_45_49351 = net_49351;
  assign seg_12_3_sp4_v_b_10_45257 = seg_12_1_sp4_v_b_34_45257;
  assign seg_12_3_sp4_v_b_11_45258 = seg_12_2_sp4_v_b_22_45258;
  assign seg_12_3_sp4_v_b_12_45259 = net_45259;
  assign seg_12_3_sp4_v_b_24_45389 = net_45389;
  assign seg_12_3_sp4_v_b_30_45395 = net_45395;
  assign seg_12_3_sp4_v_b_40_45515 = net_45515;
  assign seg_12_4_lutff_0_out_45487 = net_45487;
  assign seg_12_4_lutff_3_out_45490 = net_45490;
  assign seg_12_4_lutff_4_out_45491 = net_45491;
  assign seg_12_4_lutff_5_out_45492 = net_45492;
  assign seg_12_4_neigh_op_bot_4_45368 = seg_12_3_lutff_4_out_45368;
  assign seg_12_4_neigh_op_bot_6_45370 = seg_12_3_lutff_6_out_45370;
  assign seg_12_4_neigh_op_rgt_0_49318 = seg_13_4_lutff_0_out_49318;
  assign seg_12_4_neigh_op_rgt_3_49321 = seg_13_4_lutff_3_out_49321;
  assign seg_12_4_neigh_op_tnl_3_41782 = seg_11_5_lutff_3_out_41782;
  assign seg_12_4_sp4_h_r_11_49456 = seg_13_4_sp4_h_r_22_49456;
  assign seg_12_4_sp4_h_r_14_45627 = net_45627;
  assign seg_12_4_sp4_h_r_18_45631 = net_45631;
  assign seg_12_4_sp4_h_r_34_41793 = seg_10_4_sp4_h_r_10_41793;
  assign seg_12_4_sp4_h_r_5_49460 = seg_13_4_sp4_h_r_16_49460;
  assign seg_12_4_sp4_h_r_6_49461 = seg_14_4_sp4_h_r_30_49461;
  assign seg_12_4_sp4_h_r_9_49464 = seg_13_4_sp4_h_r_20_49464;
  assign seg_12_4_sp4_r_v_b_29_49346 = net_49346;
  assign seg_12_4_sp4_r_v_b_4_49096 = seg_12_1_sp4_r_v_b_41_49096;
  assign seg_12_4_sp4_v_b_10_45271 = seg_12_2_sp4_v_b_34_45271;
  assign seg_12_4_sp4_v_b_1_45259 = seg_12_3_sp4_v_b_12_45259;
  assign seg_12_4_sp4_v_b_36_45634 = net_45634;
  assign seg_12_4_sp4_v_t_46_45767 = seg_11_6_sp4_r_v_b_35_45767;
  assign seg_12_5_neigh_op_bnr_4_49322 = seg_13_4_lutff_4_out_49322;
  assign seg_12_5_sp4_h_r_0_49576 = net_49576;
  assign seg_12_5_sp4_h_r_10_49578 = net_49578;
  assign seg_12_5_sp4_r_v_b_13_49343 = net_49343;
  assign seg_12_5_sp4_r_v_b_21_49351 = seg_12_3_sp4_r_v_b_45_49351;
  assign seg_12_5_sp4_v_b_0_45389 = seg_12_3_sp4_v_b_24_45389;
  assign seg_12_5_sp4_v_b_36_45757 = net_45757;
  assign seg_12_5_sp4_v_b_3_45390 = seg_12_2_sp4_v_b_38_45390;
  assign seg_12_5_sp4_v_b_5_45392 = seg_12_2_sp4_v_b_40_45392;
  assign seg_12_5_sp4_v_b_6_45395 = seg_12_3_sp4_v_b_30_45395;
  assign seg_12_5_sp4_v_t_41_45885 = seg_11_8_sp4_r_v_b_17_45885;
  assign seg_12_5_sp4_v_t_45_45889 = seg_11_8_sp4_r_v_b_21_45889;
  assign seg_12_6_lutff_0_out_45733 = net_45733;
  assign seg_12_6_lutff_1_out_45734 = net_45734;
  assign seg_12_6_lutff_2_out_45735 = net_45735;
  assign seg_12_6_lutff_3_out_45736 = net_45736;
  assign seg_12_6_lutff_7_out_45740 = net_45740;
  assign seg_12_6_sp12_v_b_12_48932 = net_48932;
  assign seg_12_6_sp12_v_t_23_49698 = seg_12_16_sp12_v_b_4_49698;
  assign seg_12_6_sp4_h_l_37_34375 = seg_10_6_sp4_h_r_24_34375;
  assign seg_12_6_sp4_h_r_20_45879 = seg_14_6_sp4_h_r_44_45879;
  assign seg_12_6_sp4_h_r_3_49704 = seg_15_6_sp4_h_r_38_49704;
  assign seg_12_6_sp4_h_r_40_38213 = net_38213;
  assign seg_12_6_sp4_h_r_7_49708 = seg_15_6_sp4_h_r_42_49708;
  assign seg_12_6_sp4_v_b_40_45884 = net_45884;
  assign seg_12_6_sp4_v_b_42_45886 = net_45886;
  assign seg_12_6_sp4_v_b_44_45888 = net_45888;
  assign seg_12_6_sp4_v_b_5_45515 = seg_12_3_sp4_v_b_40_45515;
  assign seg_12_6_sp4_v_t_41_46008 = seg_11_7_sp4_r_v_b_41_46008;
  assign seg_12_6_sp4_v_t_44_46011 = seg_11_8_sp4_r_v_b_33_46011;
  assign seg_12_7_lutff_0_out_45856 = net_45856;
  assign seg_12_7_lutff_1_out_45857 = net_45857;
  assign seg_12_7_lutff_6_out_45862 = net_45862;
  assign seg_12_7_lutff_7_out_45863 = net_45863;
  assign seg_12_7_neigh_op_tnl_0_42148 = seg_11_8_lutff_0_out_42148;
  assign seg_12_7_sp4_h_r_22_45994 = net_45994;
  assign seg_12_7_sp4_h_r_24_42160 = net_42160;
  assign seg_12_7_sp4_h_r_40_38336 = seg_10_7_sp4_h_r_16_38336;
  assign seg_12_7_sp4_h_r_4_49828 = seg_14_7_sp4_h_r_28_49828;
  assign seg_12_7_sp4_r_v_b_5_49469 = seg_13_4_sp4_v_b_40_49469;
  assign seg_12_7_sp4_v_b_19_45764 = seg_11_5_sp4_r_v_b_43_45764;
  assign seg_12_7_sp4_v_b_1_45634 = seg_12_4_sp4_v_b_36_45634;
  assign seg_12_8_neigh_op_lft_0_42148 = seg_11_8_lutff_0_out_42148;
  assign seg_12_8_neigh_op_lft_2_42150 = seg_11_8_lutff_2_out_42150;
  assign seg_12_8_sp4_h_r_0_49945 = net_49945;
  assign seg_12_8_sp4_h_r_5_49952 = seg_15_8_sp4_h_r_40_49952;
  assign seg_12_8_sp4_h_r_8_49955 = net_49955;
  assign seg_12_8_sp4_h_r_9_49956 = seg_13_8_sp4_h_r_20_49956;
  assign seg_12_8_sp4_r_v_b_27_49836 = net_49836;
  assign seg_12_8_sp4_v_b_1_45757 = seg_12_5_sp4_v_b_36_45757;
  assign seg_12_8_sp4_v_b_46_46136 = net_46136;
  assign seg_12_8_sp4_v_b_6_45764 = seg_11_5_sp4_r_v_b_43_45764;
  assign seg_12_8_sp4_v_t_36_46249 = seg_11_12_sp4_r_v_b_1_46249;
  assign seg_12_9_sp4_h_r_28_42412 = net_42412;
  assign seg_12_9_sp4_h_r_32_42416 = net_42416;
  assign seg_12_9_sp4_r_v_b_43_50087 = net_50087;
  assign seg_12_9_sp4_v_b_5_45884 = seg_12_6_sp4_v_b_40_45884;
  assign seg_12_9_sp4_v_b_7_45886 = seg_12_6_sp4_v_b_42_45886;
  assign seg_12_9_sp4_v_b_9_45888 = seg_12_6_sp4_v_b_44_45888;
  assign seg_13_0_span4_vert_20_49073 = net_49073;
  assign seg_13_0_span4_vert_4_49094 = net_49094;
  assign seg_13_10_lutff_1_out_50057 = net_50057;
  assign seg_13_10_lutff_2_out_50058 = net_50058;
  assign seg_13_10_lutff_5_out_50061 = net_50061;
  assign seg_13_10_sp12_v_b_16_53529 = net_53529;
  assign seg_13_10_sp4_r_v_b_25_53911 = net_53911;
  assign seg_13_10_sp4_r_v_b_6_53672 = seg_13_7_sp4_r_v_b_43_53672;
  assign seg_13_10_sp4_r_v_b_9_53673 = seg_14_7_sp4_v_b_44_53673;
  assign seg_13_10_sp4_v_b_40_50207 = seg_12_13_sp4_r_v_b_5_50207;
  assign seg_13_10_sp4_v_b_6_49841 = seg_13_8_sp4_v_b_30_49841;
  assign seg_13_11_neigh_op_bot_5_50061 = seg_13_10_lutff_5_out_50061;
  assign seg_13_11_neigh_op_top_4_50306 = seg_13_12_lutff_4_out_50306;
  assign seg_13_11_sp12_v_b_18_53774 = net_53774;
  assign seg_13_11_sp12_v_b_20_53898 = net_53898;
  assign seg_13_11_sp4_h_r_4_54151 = seg_15_11_sp4_h_r_28_54151;
  assign seg_13_11_sp4_h_r_8_54155 = net_54155;
  assign seg_13_11_sp4_r_v_b_11_53798 = seg_14_8_sp4_v_b_46_53798;
  assign seg_13_11_sp4_v_b_10_49968 = net_49968;
  assign seg_13_11_sp4_v_b_29_50207 = seg_12_13_sp4_r_v_b_5_50207;
  assign seg_13_11_sp4_v_b_44_50334 = net_50334;
  assign seg_13_11_sp4_v_t_37_50450 = seg_12_14_sp4_r_v_b_13_50450;
  assign seg_13_11_sp4_v_t_38_50451 = seg_12_15_sp4_r_v_b_3_50451;
  assign seg_13_11_sp4_v_t_40_50453 = seg_12_15_sp4_r_v_b_5_50453;
  assign seg_13_11_sp4_v_t_42_50455 = seg_12_15_sp4_r_v_b_7_50455;
  assign seg_13_12_lutff_0_out_50302 = net_50302;
  assign seg_13_12_lutff_2_out_50304 = net_50304;
  assign seg_13_12_lutff_3_out_50305 = net_50305;
  assign seg_13_12_lutff_4_out_50306 = net_50306;
  assign seg_13_12_lutff_5_out_50307 = net_50307;
  assign seg_13_12_lutff_6_out_50308 = net_50308;
  assign seg_13_12_sp12_v_b_1_52762 = seg_13_1_sp12_v_b_22_52762;
  assign seg_13_12_sp4_h_r_34_46608 = net_46608;
  assign seg_13_12_sp4_r_v_b_31_54163 = net_54163;
  assign seg_13_12_sp4_v_b_10_50091 = seg_12_11_sp4_r_v_b_23_50091;
  assign seg_13_12_sp4_v_b_7_50086 = seg_12_10_sp4_r_v_b_31_50086;
  assign seg_13_12_sp4_v_t_37_50573 = seg_12_13_sp4_r_v_b_37_50573;
  assign seg_13_12_sp4_v_t_39_50575 = seg_12_15_sp4_r_v_b_15_50575;
  assign seg_13_12_sp4_v_t_45_50581 = seg_12_15_sp4_r_v_b_21_50581;
  assign seg_13_13_lutff_0_out_50425 = net_50425;
  assign seg_13_13_lutff_2_out_50427 = net_50427;
  assign seg_13_13_lutff_3_out_50428 = net_50428;
  assign seg_13_13_lutff_5_out_50430 = net_50430;
  assign seg_13_13_neigh_op_bot_0_50302 = seg_13_12_lutff_0_out_50302;
  assign seg_13_13_neigh_op_bot_2_50304 = seg_13_12_lutff_2_out_50304;
  assign seg_13_13_neigh_op_bot_3_50305 = seg_13_12_lutff_3_out_50305;
  assign seg_13_13_neigh_op_bot_6_50308 = seg_13_12_lutff_6_out_50308;
  assign seg_13_13_neigh_op_lft_2_46596 = seg_12_13_lutff_2_out_46596;
  assign seg_13_13_sp4_h_r_3_54396 = seg_14_13_sp4_h_r_14_54396;
  assign seg_13_13_sp4_r_v_b_31_54286 = net_54286;
  assign seg_13_13_sp4_r_v_b_41_54408 = net_54408;
  assign seg_13_13_sp4_v_b_10_50214 = seg_12_10_sp4_r_v_b_47_50214;
  assign seg_13_13_sp4_v_b_2_50206 = seg_12_10_sp4_r_v_b_39_50206;
  assign seg_13_13_sp4_v_b_34_50460 = net_50460;
  assign seg_13_13_sp4_v_b_44_50580 = net_50580;
  assign seg_13_13_sp4_v_b_5_50207 = seg_12_13_sp4_r_v_b_5_50207;
  assign seg_13_13_sp4_v_b_8_50212 = seg_12_10_sp4_r_v_b_45_50212;
  assign seg_13_13_sp4_v_t_42_50701 = seg_12_15_sp4_r_v_b_31_50701;
  assign seg_13_14_lutff_1_out_50549 = net_50549;
  assign seg_13_14_lutff_2_out_50550 = net_50550;
  assign seg_13_14_neigh_op_bnl_2_46596 = seg_12_13_lutff_2_out_46596;
  assign seg_13_14_neigh_op_tnl_0_46840 = seg_12_15_lutff_0_out_46840;
  assign seg_13_14_neigh_op_tnr_2_54504 = seg_14_15_lutff_2_out_54504;
  assign seg_13_14_sp12_v_b_10_53651 = net_53651;
  assign seg_13_14_sp12_v_b_14_53897 = net_53897;
  assign seg_13_14_sp4_h_r_0_54514 = seg_15_14_sp4_h_r_24_54514;
  assign seg_13_14_sp4_h_r_10_54516 = seg_15_14_sp4_h_r_34_54516;
  assign seg_13_14_sp4_h_r_18_50692 = net_50692;
  assign seg_13_14_sp4_h_r_28_46858 = net_46858;
  assign seg_13_14_sp4_h_r_2_54518 = net_54518;
  assign seg_13_14_sp4_h_r_34_46854 = net_46854;
  assign seg_13_14_sp4_h_r_40_43028 = net_43028;
  assign seg_13_14_sp4_h_r_4_54520 = seg_15_14_sp4_h_r_28_54520;
  assign seg_13_14_sp4_r_v_b_35_54413 = net_54413;
  assign seg_13_14_sp4_r_v_b_3_54159 = net_54159;
  assign seg_13_14_sp4_r_v_b_7_54163 = seg_13_12_sp4_r_v_b_31_54163;
  assign seg_13_14_sp4_v_b_0_50327 = net_50327;
  assign seg_13_14_sp4_v_b_38_50697 = net_50697;
  assign seg_13_14_sp4_v_b_4_50331 = seg_12_11_sp4_r_v_b_41_50331;
  assign seg_13_14_sp4_v_b_6_50333 = seg_12_11_sp4_r_v_b_43_50333;
  assign seg_13_14_sp4_v_b_8_50335 = seg_12_11_sp4_r_v_b_45_50335;
  assign seg_13_14_sp4_v_b_9_50334 = seg_13_11_sp4_v_b_44_50334;
  assign seg_13_14_sp4_v_t_38_50820 = seg_13_17_sp4_v_b_14_50820;
  assign seg_13_15_lutff_1_out_50672 = net_50672;
  assign seg_13_15_lutff_2_out_50673 = net_50673;
  assign seg_13_15_neigh_op_bot_1_50549 = seg_13_14_lutff_1_out_50549;
  assign seg_13_15_neigh_op_lft_3_46843 = seg_12_15_lutff_3_out_46843;
  assign seg_13_15_neigh_op_lft_4_46844 = seg_12_15_lutff_4_out_46844;
  assign seg_13_15_neigh_op_rgt_2_54504 = seg_14_15_lutff_2_out_54504;
  assign seg_13_15_neigh_op_top_1_50795 = seg_13_16_lutff_1_out_50795;
  assign seg_13_15_neigh_op_top_3_50797 = seg_13_16_lutff_3_out_50797;
  assign seg_13_15_neigh_op_top_6_50800 = seg_13_16_lutff_6_out_50800;
  assign seg_13_15_sp12_v_b_16_54144 = net_54144;
  assign seg_13_15_sp4_h_l_36_39314 = seg_12_15_sp4_h_r_36_39314;
  assign seg_13_15_sp4_r_v_b_41_54654 = net_54654;
  assign seg_13_15_sp4_r_v_b_43_54656 = net_54656;
  assign seg_13_15_sp4_r_v_b_45_54658 = net_54658;
  assign seg_13_15_sp4_v_b_10_50460 = seg_13_13_sp4_v_b_34_50460;
  assign seg_13_15_sp4_v_b_13_50573 = seg_12_13_sp4_r_v_b_37_50573;
  assign seg_13_15_sp4_v_b_18_50578 = net_50578;
  assign seg_13_15_sp4_v_b_39_50821 = seg_12_17_sp4_r_v_b_15_50821;
  assign seg_13_15_sp4_v_b_46_50828 = net_50828;
  assign seg_13_15_sp4_v_t_43_50948 = seg_13_17_sp4_v_b_30_50948;
  assign seg_13_16_lutff_1_out_50795 = net_50795;
  assign seg_13_16_lutff_2_out_50796 = net_50796;
  assign seg_13_16_lutff_3_out_50797 = net_50797;
  assign seg_13_16_lutff_4_out_50798 = net_50798;
  assign seg_13_16_lutff_5_out_50799 = net_50799;
  assign seg_13_16_lutff_6_out_50800 = net_50800;
  assign seg_13_16_lutff_7_out_50801 = net_50801;
  assign seg_13_16_neigh_op_bot_1_50672 = seg_13_15_lutff_1_out_50672;
  assign seg_13_16_neigh_op_bot_2_50673 = seg_13_15_lutff_2_out_50673;
  assign seg_13_16_neigh_op_lft_4_46967 = seg_12_16_lutff_4_out_46967;
  assign seg_13_16_neigh_op_tnl_6_47092 = seg_12_17_lutff_6_out_47092;
  assign seg_13_16_neigh_op_top_3_50920 = seg_13_17_lutff_3_out_50920;
  assign seg_13_16_neigh_op_top_4_50921 = seg_13_17_lutff_4_out_50921;
  assign seg_13_16_neigh_op_top_5_50922 = seg_13_17_lutff_5_out_50922;
  assign seg_13_16_sp4_h_r_22_50932 = net_50932;
  assign seg_13_16_sp4_h_r_38_43272 = net_43272;
  assign seg_13_16_sp4_r_v_b_39_54775 = net_54775;
  assign seg_13_16_sp4_r_v_b_7_54409 = net_54409;
  assign seg_13_16_sp4_r_v_b_9_54411 = net_54411;
  assign seg_13_16_sp4_v_b_10_50583 = seg_12_15_sp4_r_v_b_23_50583;
  assign seg_13_16_sp4_v_b_38_50943 = net_50943;
  assign seg_13_16_sp4_v_b_6_50579 = seg_12_13_sp4_r_v_b_43_50579;
  assign seg_13_16_sp4_v_b_9_50580 = seg_13_13_sp4_v_b_44_50580;
  assign seg_13_16_sp4_v_t_38_51066 = seg_13_19_sp4_v_b_14_51066;
  assign seg_13_16_sp4_v_t_39_51067 = seg_13_18_sp4_v_b_26_51067;
  assign seg_13_16_sp4_v_t_45_51073 = seg_13_18_sp4_v_b_32_51073;
  assign seg_13_17_lutff_1_out_50918 = net_50918;
  assign seg_13_17_lutff_3_out_50920 = net_50920;
  assign seg_13_17_lutff_4_out_50921 = net_50921;
  assign seg_13_17_lutff_5_out_50922 = net_50922;
  assign seg_13_17_lutff_7_out_50924 = net_50924;
  assign seg_13_17_neigh_op_bot_3_50797 = seg_13_16_lutff_3_out_50797;
  assign seg_13_17_neigh_op_lft_6_47092 = seg_12_17_lutff_6_out_47092;
  assign seg_13_17_neigh_op_lft_7_47093 = seg_12_17_lutff_7_out_47093;
  assign seg_13_17_sp4_h_r_14_51057 = net_51057;
  assign seg_13_17_sp4_h_r_30_47229 = net_47229;
  assign seg_13_17_sp4_h_r_46_43393 = net_43393;
  assign seg_13_17_sp4_r_v_b_15_54652 = net_54652;
  assign seg_13_17_sp4_v_b_14_50820 = net_50820;
  assign seg_13_17_sp4_v_b_30_50948 = net_50948;
  assign seg_13_17_sp4_v_b_3_50697 = seg_13_14_sp4_v_b_38_50697;
  assign seg_13_17_sp4_v_b_7_50701 = seg_12_15_sp4_r_v_b_31_50701;
  assign seg_13_18_lutff_1_out_51041 = net_51041;
  assign seg_13_18_lutff_2_out_51042 = net_51042;
  assign seg_13_18_lutff_6_out_51046 = net_51046;
  assign seg_13_18_neigh_op_bot_7_50924 = seg_13_17_lutff_7_out_50924;
  assign seg_13_18_sp12_v_b_0_53529 = seg_13_10_sp12_v_b_16_53529;
  assign seg_13_18_sp12_v_b_2_53651 = seg_13_14_sp12_v_b_10_53651;
  assign seg_13_18_sp12_v_b_5_53774 = seg_13_11_sp12_v_b_18_53774;
  assign seg_13_18_sp12_v_b_6_53897 = seg_13_14_sp12_v_b_14_53897;
  assign seg_13_18_sp12_v_b_7_53898 = seg_13_11_sp12_v_b_20_53898;
  assign seg_13_18_sp4_h_r_14_51180 = net_51180;
  assign seg_13_18_sp4_h_r_38_43518 = net_43518;
  assign seg_13_18_sp4_r_v_b_4_54654 = seg_13_15_sp4_r_v_b_41_54654;
  assign seg_13_18_sp4_r_v_b_6_54656 = seg_13_15_sp4_r_v_b_43_54656;
  assign seg_13_18_sp4_r_v_b_8_54658 = seg_13_15_sp4_r_v_b_45_54658;
  assign seg_13_18_sp4_v_b_11_50828 = seg_13_15_sp4_v_b_46_50828;
  assign seg_13_18_sp4_v_b_26_51067 = net_51067;
  assign seg_13_18_sp4_v_b_32_51073 = net_51073;
  assign seg_13_18_sp4_v_b_3_50820 = seg_13_17_sp4_v_b_14_50820;
  assign seg_13_19_sp4_v_b_14_51066 = net_51066;
  assign seg_13_19_sp4_v_b_3_50943 = seg_13_16_sp4_v_b_38_50943;
  assign seg_13_19_sp4_v_b_6_50948 = seg_13_17_sp4_v_b_30_50948;
  assign seg_13_1_lutff_3_out_48911 = net_48911;
  assign seg_13_1_lutff_5_out_48913 = net_48913;
  assign seg_13_1_neigh_op_top_2_49038 = seg_13_2_lutff_2_out_49038;
  assign seg_13_1_neigh_op_top_3_49039 = seg_13_2_lutff_3_out_49039;
  assign seg_13_1_neigh_op_top_4_49040 = seg_13_2_lutff_4_out_49040;
  assign seg_13_1_sp12_v_b_22_52762 = net_52762;
  assign seg_13_1_sp4_h_r_22_49051 = net_49051;
  assign seg_13_1_sp4_h_r_44_41397 = net_41397;
  assign seg_13_1_sp4_v_b_38_49092 = net_49092;
  assign seg_13_1_sp4_v_b_4_49094 = seg_13_0_span4_vert_4_49094;
  assign seg_13_23_sp12_v_b_0_54144 = seg_13_15_sp12_v_b_16_54144;
  assign seg_13_2_lutff_0_out_49036 = net_49036;
  assign seg_13_2_lutff_1_out_49037 = net_49037;
  assign seg_13_2_lutff_2_out_49038 = net_49038;
  assign seg_13_2_lutff_3_out_49039 = net_49039;
  assign seg_13_2_lutff_4_out_49040 = net_49040;
  assign seg_13_2_neigh_op_bnl_2_45079 = seg_12_1_lutff_2_out_45079;
  assign seg_13_2_neigh_op_bnl_3_45080 = seg_12_1_lutff_3_out_45080;
  assign seg_13_2_neigh_op_bot_3_48911 = seg_13_1_lutff_3_out_48911;
  assign seg_13_2_neigh_op_top_7_49202 = seg_13_3_lutff_7_out_49202;
  assign seg_13_2_sp4_h_l_41_37720 = seg_11_2_sp4_h_r_28_37720;
  assign seg_13_2_sp4_h_l_47_37716 = seg_11_2_sp4_h_r_34_37716;
  assign seg_13_2_sp4_r_v_b_25_52921 = net_52921;
  assign seg_13_2_sp4_r_v_b_37_53051 = net_53051;
  assign seg_13_2_sp4_v_b_10_49076 = seg_12_1_sp4_r_v_b_23_49076;
  assign seg_13_2_sp4_v_b_6_49071 = seg_12_1_sp4_r_v_b_19_49071;
  assign seg_13_2_sp4_v_b_8_49074 = seg_12_1_sp4_r_v_b_21_49074;
  assign seg_13_2_sp4_v_b_9_49073 = seg_13_0_span4_vert_20_49073;
  assign seg_13_3_lutff_0_out_49195 = net_49195;
  assign seg_13_3_lutff_1_out_49196 = net_49196;
  assign seg_13_3_lutff_2_out_49197 = net_49197;
  assign seg_13_3_lutff_4_out_49199 = net_49199;
  assign seg_13_3_lutff_6_out_49201 = net_49201;
  assign seg_13_3_lutff_7_out_49202 = net_49202;
  assign seg_13_3_neigh_op_tnl_5_45492 = seg_12_4_lutff_5_out_45492;
  assign seg_13_3_neigh_op_tnr_2_53151 = seg_14_4_lutff_2_out_53151;
  assign seg_13_3_sp4_h_r_10_53163 = net_53163;
  assign seg_13_3_sp4_h_r_16_49337 = seg_15_3_sp4_h_r_40_49337;
  assign seg_13_3_sp4_h_r_1_53162 = seg_16_3_sp4_h_r_36_53162;
  assign seg_13_3_sp4_h_r_2_53165 = net_53165;
  assign seg_13_3_sp4_r_v_b_35_53060 = net_53060;
  assign seg_13_3_sp4_v_b_11_49089 = seg_12_1_sp4_r_v_b_35_49089;
  assign seg_13_3_sp4_v_b_17_49096 = seg_12_1_sp4_r_v_b_41_49096;
  assign seg_13_3_sp4_v_b_1_49078 = seg_12_1_sp4_r_v_b_25_49078;
  assign seg_13_3_sp4_v_b_34_49230 = net_49230;
  assign seg_13_3_sp4_v_t_38_49467 = seg_13_4_sp4_v_b_38_49467;
  assign seg_13_4_lutff_0_out_49318 = net_49318;
  assign seg_13_4_lutff_3_out_49321 = net_49321;
  assign seg_13_4_lutff_4_out_49322 = net_49322;
  assign seg_13_4_lutff_5_out_49323 = net_49323;
  assign seg_13_4_lutff_6_out_49324 = net_49324;
  assign seg_13_4_sp12_h_r_10_34126 = seg_11_4_sp12_h_r_6_34126;
  assign seg_13_4_sp4_h_l_41_37966 = seg_11_4_sp4_h_r_28_37966;
  assign seg_13_4_sp4_h_r_16_49460 = net_49460;
  assign seg_13_4_sp4_h_r_20_49464 = net_49464;
  assign seg_13_4_sp4_h_r_22_49456 = net_49456;
  assign seg_13_4_sp4_h_r_32_45632 = seg_11_4_sp4_h_r_8_45632;
  assign seg_13_4_sp4_h_r_36_41792 = net_41792;
  assign seg_13_4_sp4_h_r_38_41796 = net_41796;
  assign seg_13_4_sp4_h_r_4_53290 = net_53290;
  assign seg_13_4_sp4_h_r_8_53294 = net_53294;
  assign seg_13_4_sp4_h_r_9_53295 = seg_14_4_sp4_h_r_20_53295;
  assign seg_13_4_sp4_r_v_b_13_53051 = seg_13_2_sp4_r_v_b_37_53051;
  assign seg_13_4_sp4_r_v_b_15_53053 = net_53053;
  assign seg_13_4_sp4_r_v_b_1_52921 = seg_13_2_sp4_r_v_b_25_52921;
  assign seg_13_4_sp4_r_v_b_35_53183 = net_53183;
  assign seg_13_4_sp4_r_v_b_41_53301 = net_53301;
  assign seg_13_4_sp4_v_b_0_49091 = seg_12_1_sp4_r_v_b_37_49091;
  assign seg_13_4_sp4_v_b_1_49090 = seg_12_2_sp4_r_v_b_25_49090;
  assign seg_13_4_sp4_v_b_2_49093 = seg_12_1_sp4_r_v_b_39_49093;
  assign seg_13_4_sp4_v_b_38_49467 = net_49467;
  assign seg_13_4_sp4_v_b_3_49092 = seg_13_1_sp4_v_b_38_49092;
  assign seg_13_4_sp4_v_b_40_49469 = net_49469;
  assign seg_13_4_sp4_v_b_4_49096 = seg_12_1_sp4_r_v_b_41_49096;
  assign seg_13_5_lutff_0_out_49441 = net_49441;
  assign seg_13_5_lutff_1_out_49442 = net_49442;
  assign seg_13_5_neigh_op_bot_3_49321 = seg_13_4_lutff_3_out_49321;
  assign seg_13_5_sp4_h_l_39_38087 = seg_11_5_sp4_h_r_26_38087;
  assign seg_13_5_sp4_h_r_34_45747 = seg_11_5_sp4_h_r_10_45747;
  assign seg_13_5_sp4_r_v_b_45_53428 = net_53428;
  assign seg_13_5_sp4_v_b_10_49230 = seg_13_3_sp4_v_b_34_49230;
  assign seg_13_5_sp4_v_b_1_49219 = seg_12_3_sp4_r_v_b_25_49219;
  assign seg_13_5_sp4_v_b_26_49468 = net_49468;
  assign seg_13_5_sp4_v_b_4_49224 = seg_12_2_sp4_r_v_b_41_49224;
  assign seg_13_6_neigh_op_bot_1_49442 = seg_13_5_lutff_1_out_49442;
  assign seg_13_6_neigh_op_tnl_1_45857 = seg_12_7_lutff_1_out_45857;
  assign seg_13_6_sp4_h_r_0_53530 = net_53530;
  assign seg_13_6_sp4_h_r_10_53532 = net_53532;
  assign seg_13_6_sp4_h_r_20_49710 = net_49710;
  assign seg_13_6_sp4_h_r_26_45872 = seg_11_6_sp4_h_r_2_45872;
  assign seg_13_6_sp4_h_r_2_53534 = net_53534;
  assign seg_13_6_sp4_h_r_30_45876 = net_45876;
  assign seg_13_6_sp4_h_r_44_42048 = net_42048;
  assign seg_13_6_sp4_h_r_8_53540 = net_53540;
  assign seg_13_6_sp4_r_v_b_7_53179 = net_53179;
  assign seg_13_6_sp4_v_b_0_49343 = seg_12_5_sp4_r_v_b_13_49343;
  assign seg_13_6_sp4_v_b_5_49346 = seg_12_4_sp4_r_v_b_29_49346;
  assign seg_13_6_sp4_v_t_38_49836 = seg_12_8_sp4_r_v_b_27_49836;
  assign seg_13_7_lutff_0_out_49687 = net_49687;
  assign seg_13_7_lutff_3_out_49690 = net_49690;
  assign seg_13_7_lutff_6_out_49693 = net_49693;
  assign seg_13_7_neigh_op_lft_0_45856 = seg_12_7_lutff_0_out_45856;
  assign seg_13_7_neigh_op_lft_7_45863 = seg_12_7_lutff_7_out_45863;
  assign seg_13_7_neigh_op_rgt_6_53524 = seg_14_7_lutff_6_out_53524;
  assign seg_13_7_sp4_h_l_40_38336 = seg_10_7_sp4_h_r_16_38336;
  assign seg_13_7_sp4_h_r_14_49827 = net_49827;
  assign seg_13_7_sp4_h_r_1_53654 = seg_14_7_sp4_h_r_12_53654;
  assign seg_13_7_sp4_h_r_2_53657 = net_53657;
  assign seg_13_7_sp4_r_v_b_21_53428 = seg_13_5_sp4_r_v_b_45_53428;
  assign seg_13_7_sp4_r_v_b_37_53666 = net_53666;
  assign seg_13_7_sp4_r_v_b_41_53670 = net_53670;
  assign seg_13_7_sp4_r_v_b_43_53672 = net_53672;
  assign seg_13_7_sp4_v_b_2_49468 = seg_13_5_sp4_v_b_26_49468;
  assign seg_13_7_sp4_v_b_3_49467 = seg_13_4_sp4_v_b_38_49467;
  assign seg_13_8_lutff_5_out_49815 = net_49815;
  assign seg_13_8_lutff_6_out_49816 = net_49816;
  assign seg_13_8_neigh_op_bot_3_49690 = seg_13_7_lutff_3_out_49690;
  assign seg_13_8_neigh_op_bot_6_49693 = seg_13_7_lutff_6_out_49693;
  assign seg_13_8_neigh_op_top_2_49935 = seg_13_9_lutff_2_out_49935;
  assign seg_13_8_neigh_op_top_5_49938 = seg_13_9_lutff_5_out_49938;
  assign seg_13_8_sp4_h_l_38_38457 = seg_10_8_sp4_h_r_14_38457;
  assign seg_13_8_sp4_h_r_0_53776 = seg_15_8_sp4_h_r_24_53776;
  assign seg_13_8_sp4_h_r_11_53779 = seg_14_8_sp4_h_r_22_53779;
  assign seg_13_8_sp4_h_r_20_49956 = net_49956;
  assign seg_13_8_sp4_h_r_24_46114 = net_46114;
  assign seg_13_8_sp4_h_r_2_53780 = net_53780;
  assign seg_13_8_sp4_h_r_32_46124 = net_46124;
  assign seg_13_8_sp4_v_b_30_49841 = net_49841;
  assign seg_13_8_sp4_v_t_43_50087 = seg_12_9_sp4_r_v_b_43_50087;
  assign seg_13_9_lutff_2_out_49935 = net_49935;
  assign seg_13_9_lutff_5_out_49938 = net_49938;
  assign seg_13_9_sp4_h_r_11_53902 = seg_16_9_sp4_h_r_46_53902;
  assign seg_13_9_sp4_h_r_7_53908 = seg_16_9_sp4_h_r_42_53908;
  assign seg_13_9_sp4_v_t_40_50207 = seg_12_13_sp4_r_v_b_5_50207;
  assign seg_14_0_span4_horz_r_0_56601 = seg_17_0_span4_horz_r_12_56601;
  assign seg_14_10_sp12_h_r_2_54019 = net_54019;
  assign seg_14_10_sp4_h_r_14_54027 = net_54027;
  assign seg_14_10_sp4_h_r_16_54029 = net_54029;
  assign seg_14_10_sp4_h_r_18_54031 = net_54031;
  assign seg_14_10_sp4_h_r_20_54033 = net_54033;
  assign seg_14_10_sp4_h_r_22_54025 = net_54025;
  assign seg_14_10_sp4_r_v_b_13_57619 = net_57619;
  assign seg_14_10_sp4_r_v_b_27_57743 = net_57743;
  assign seg_14_10_sp4_r_v_b_29_57745 = net_57745;
  assign seg_14_10_sp4_r_v_b_31_57747 = net_57747;
  assign seg_14_10_sp4_r_v_b_35_57751 = net_57751;
  assign seg_14_10_sp4_v_b_0_53666 = seg_13_7_sp4_r_v_b_37_53666;
  assign seg_14_10_sp4_v_b_32_53920 = seg_14_12_sp4_v_b_8_53920;
  assign seg_14_10_sp4_v_b_8_53674 = net_53674;
  assign seg_14_10_sp4_v_t_38_54159 = seg_13_14_sp4_r_v_b_3_54159;
  assign seg_14_11_sp4_h_l_40_42659 = seg_11_11_sp4_h_r_16_42659;
  assign seg_14_11_sp4_h_r_24_50314 = net_50314;
  assign seg_14_11_sp4_h_r_5_57982 = seg_15_11_sp4_h_r_16_57982;
  assign seg_14_11_sp4_r_v_b_15_57744 = net_57744;
  assign seg_14_11_sp4_r_v_b_17_57746 = net_57746;
  assign seg_14_11_sp4_r_v_b_1_57618 = seg_15_8_sp4_v_b_36_57618;
  assign seg_14_11_sp4_r_v_b_23_57752 = net_57752;
  assign seg_14_11_sp4_v_b_1_53788 = seg_14_8_sp4_v_b_36_53788;
  assign seg_14_12_lutff_4_out_54137 = net_54137;
  assign seg_14_12_neigh_op_bnr_0_57840 = seg_15_11_lutff_0_out_57840;
  assign seg_14_12_sp4_h_r_6_58106 = seg_16_12_sp4_h_r_30_58106;
  assign seg_14_12_sp4_v_b_1_53911 = seg_13_10_sp4_r_v_b_25_53911;
  assign seg_14_12_sp4_v_b_40_54284 = net_54284;
  assign seg_14_12_sp4_v_b_8_53920 = net_53920;
  assign seg_14_12_sp4_v_t_42_54409 = seg_13_16_sp4_r_v_b_7_54409;
  assign seg_14_13_lutff_0_out_54256 = net_54256;
  assign seg_14_13_lutff_1_out_54257 = net_54257;
  assign seg_14_13_lutff_3_out_54259 = net_54259;
  assign seg_14_13_lutff_4_out_54260 = net_54260;
  assign seg_14_13_lutff_6_out_54262 = net_54262;
  assign seg_14_13_neigh_op_bot_4_54137 = seg_14_12_lutff_4_out_54137;
  assign seg_14_13_neigh_op_tnr_4_58213 = seg_15_14_lutff_4_out_58213;
  assign seg_14_13_sp12_h_r_12_35232 = net_35232;
  assign seg_14_13_sp12_v_b_12_57482 = net_57482;
  assign seg_14_13_sp4_h_r_0_58221 = net_58221;
  assign seg_14_13_sp4_h_r_10_58223 = net_58223;
  assign seg_14_13_sp4_h_r_14_54396 = net_54396;
  assign seg_14_13_sp4_h_r_36_46730 = net_46730;
  assign seg_14_13_sp4_h_r_46_46732 = net_46732;
  assign seg_14_13_sp4_r_v_b_21_57996 = net_57996;
  assign seg_14_13_sp4_r_v_b_29_58114 = net_58114;
  assign seg_14_13_sp4_r_v_b_31_58116 = net_58116;
  assign seg_14_13_sp4_r_v_b_39_58236 = net_58236;
  assign seg_14_13_sp4_v_b_32_54289 = seg_14_15_sp4_v_b_8_54289;
  assign seg_14_13_sp4_v_b_44_54411 = seg_13_16_sp4_r_v_b_9_54411;
  assign seg_14_14_lutff_0_out_54379 = net_54379;
  assign seg_14_14_lutff_2_out_54381 = net_54381;
  assign seg_14_14_lutff_4_out_54383 = net_54383;
  assign seg_14_14_lutff_5_out_54384 = net_54384;
  assign seg_14_14_lutff_6_out_54385 = net_54385;
  assign seg_14_14_lutff_7_out_54386 = net_54386;
  assign seg_14_14_neigh_op_bot_3_54259 = seg_14_13_lutff_3_out_54259;
  assign seg_14_14_neigh_op_bot_6_54262 = seg_14_13_lutff_6_out_54262;
  assign seg_14_14_neigh_op_lft_1_50549 = seg_13_14_lutff_1_out_50549;
  assign seg_14_14_sp12_v_b_12_57605 = net_57605;
  assign seg_14_14_sp4_h_l_40_43028 = seg_13_14_sp4_h_r_40_43028;
  assign seg_14_14_sp4_h_r_10_58346 = net_58346;
  assign seg_14_14_sp4_h_r_30_50691 = net_50691;
  assign seg_14_14_sp4_h_r_4_58350 = net_58350;
  assign seg_14_14_sp4_h_r_8_58354 = net_58354;
  assign seg_14_14_sp4_r_v_b_1_57987 = net_57987;
  assign seg_14_14_sp4_r_v_b_33_58241 = net_58241;
  assign seg_14_14_sp4_r_v_b_37_58357 = net_58357;
  assign seg_14_14_sp4_r_v_b_41_58361 = net_58361;
  assign seg_14_14_sp4_r_v_b_43_58363 = net_58363;
  assign seg_14_14_sp4_r_v_b_47_58367 = net_58367;
  assign seg_14_14_sp4_v_b_16_54284 = seg_14_12_sp4_v_b_40_54284;
  assign seg_14_14_sp4_v_b_33_54411 = seg_13_16_sp4_r_v_b_9_54411;
  assign seg_14_14_sp4_v_b_3_54159 = seg_13_14_sp4_r_v_b_3_54159;
  assign seg_14_14_sp4_v_t_39_54652 = seg_13_17_sp4_r_v_b_15_54652;
  assign seg_14_15_lutff_0_out_54502 = net_54502;
  assign seg_14_15_lutff_2_out_54504 = net_54504;
  assign seg_14_15_lutff_3_out_54505 = net_54505;
  assign seg_14_15_lutff_4_out_54506 = net_54506;
  assign seg_14_15_lutff_5_out_54507 = net_54507;
  assign seg_14_15_lutff_6_out_54508 = net_54508;
  assign seg_14_15_lutff_7_out_54509 = net_54509;
  assign seg_14_15_neigh_op_bot_0_54379 = seg_14_14_lutff_0_out_54379;
  assign seg_14_15_neigh_op_bot_2_54381 = seg_14_14_lutff_2_out_54381;
  assign seg_14_15_neigh_op_bot_4_54383 = seg_14_14_lutff_4_out_54383;
  assign seg_14_15_neigh_op_bot_5_54384 = seg_14_14_lutff_5_out_54384;
  assign seg_14_15_neigh_op_bot_6_54385 = seg_14_14_lutff_6_out_54385;
  assign seg_14_15_neigh_op_bot_7_54386 = seg_14_14_lutff_7_out_54386;
  assign seg_14_15_sp12_v_b_18_58096 = net_58096;
  assign seg_14_15_sp4_h_l_43_43152 = seg_12_15_sp4_h_r_30_43152;
  assign seg_14_15_sp4_h_r_36_46976 = net_46976;
  assign seg_14_15_sp4_r_v_b_15_58236 = seg_14_13_sp4_r_v_b_39_58236;
  assign seg_14_15_sp4_r_v_b_5_58114 = seg_14_13_sp4_r_v_b_29_58114;
  assign seg_14_15_sp4_v_b_7_54286 = seg_13_13_sp4_r_v_b_31_54286;
  assign seg_14_15_sp4_v_b_8_54289 = net_54289;
  assign seg_14_15_sp4_v_t_39_54775 = seg_13_16_sp4_r_v_b_39_54775;
  assign seg_14_16_neigh_op_bot_0_54502 = seg_14_15_lutff_0_out_54502;
  assign seg_14_16_neigh_op_bot_3_54505 = seg_14_15_lutff_3_out_54505;
  assign seg_14_16_neigh_op_bot_5_54507 = seg_14_15_lutff_5_out_54507;
  assign seg_14_16_neigh_op_bot_6_54508 = seg_14_15_lutff_6_out_54508;
  assign seg_14_16_neigh_op_bot_7_54509 = seg_14_15_lutff_7_out_54509;
  assign seg_14_16_neigh_op_tnr_2_58580 = seg_15_17_lutff_2_out_58580;
  assign seg_14_16_neigh_op_top_7_54755 = seg_14_17_lutff_7_out_54755;
  assign seg_14_16_sp4_h_l_38_43272 = seg_13_16_sp4_h_r_38_43272;
  assign seg_14_16_sp4_h_r_10_58592 = seg_16_16_sp4_h_r_34_58592;
  assign seg_14_16_sp4_h_r_14_54765 = net_54765;
  assign seg_14_16_sp4_h_r_20_54771 = seg_16_16_sp4_h_r_44_54771;
  assign seg_14_16_sp4_h_r_24_50929 = net_50929;
  assign seg_14_16_sp4_h_r_4_58596 = net_58596;
  assign seg_14_16_sp4_h_r_8_58600 = seg_16_16_sp4_h_r_32_58600;
  assign seg_14_16_sp4_r_v_b_11_58243 = net_58243;
  assign seg_14_16_sp4_r_v_b_27_58481 = seg_14_18_sp4_r_v_b_3_58481;
  assign seg_14_16_sp4_r_v_b_29_58483 = seg_14_18_sp4_r_v_b_5_58483;
  assign seg_14_16_sp4_r_v_b_39_58605 = net_58605;
  assign seg_14_16_sp4_v_b_11_54413 = seg_13_14_sp4_r_v_b_35_54413;
  assign seg_14_16_sp4_v_b_34_54660 = seg_14_18_sp4_v_b_10_54660;
  assign seg_14_16_sp4_v_b_36_54772 = seg_14_18_sp4_v_b_12_54772;
  assign seg_14_16_sp4_v_b_44_54780 = net_54780;
  assign seg_14_16_sp4_v_b_4_54408 = seg_13_13_sp4_r_v_b_41_54408;
  assign seg_14_16_sp4_v_t_46_54905 = seg_14_19_sp4_v_b_22_54905;
  assign seg_14_17_lutff_2_out_54750 = net_54750;
  assign seg_14_17_lutff_3_out_54751 = net_54751;
  assign seg_14_17_lutff_5_out_54753 = net_54753;
  assign seg_14_17_lutff_6_out_54754 = net_54754;
  assign seg_14_17_lutff_7_out_54755 = net_54755;
  assign seg_14_17_neigh_op_top_1_54872 = seg_14_18_lutff_1_out_54872;
  assign seg_14_17_neigh_op_top_7_54878 = seg_14_18_lutff_7_out_54878;
  assign seg_14_17_sp4_h_r_0_58713 = net_58713;
  assign seg_14_17_sp4_h_r_11_58716 = seg_17_17_sp4_h_r_46_58716;
  assign seg_14_17_sp4_h_r_14_54888 = seg_16_17_sp4_h_r_38_54888;
  assign seg_14_17_sp4_h_r_2_58717 = net_58717;
  assign seg_14_17_sp4_r_v_b_19_58486 = net_58486;
  assign seg_14_17_sp4_r_v_b_3_58358 = net_58358;
  assign seg_14_18_lutff_0_out_54871 = net_54871;
  assign seg_14_18_lutff_1_out_54872 = net_54872;
  assign seg_14_18_lutff_3_out_54874 = net_54874;
  assign seg_14_18_lutff_5_out_54876 = net_54876;
  assign seg_14_18_lutff_7_out_54878 = net_54878;
  assign seg_14_18_neigh_op_bot_5_54753 = seg_14_17_lutff_5_out_54753;
  assign seg_14_18_neigh_op_bot_6_54754 = seg_14_17_lutff_6_out_54754;
  assign seg_14_18_neigh_op_lft_1_51041 = seg_13_18_lutff_1_out_51041;
  assign seg_14_18_neigh_op_lft_2_51042 = seg_13_18_lutff_2_out_51042;
  assign seg_14_18_neigh_op_lft_6_51046 = seg_13_18_lutff_6_out_51046;
  assign seg_14_18_sp4_h_l_37_43513 = seg_10_18_sp4_h_r_0_43513;
  assign seg_14_18_sp4_h_l_45_43523 = seg_10_18_sp4_h_r_8_43523;
  assign seg_14_18_sp4_h_r_9_58847 = seg_17_18_sp4_h_r_44_58847;
  assign seg_14_18_sp4_r_v_b_11_58489 = net_58489;
  assign seg_14_18_sp4_r_v_b_13_58603 = net_58603;
  assign seg_14_18_sp4_r_v_b_14_58604 = seg_15_16_sp4_v_b_38_58604;
  assign seg_14_18_sp4_r_v_b_15_58605 = seg_14_16_sp4_r_v_b_39_58605;
  assign seg_14_18_sp4_r_v_b_20_58610 = seg_15_16_sp4_v_b_44_58610;
  assign seg_14_18_sp4_r_v_b_3_58481 = net_58481;
  assign seg_14_18_sp4_r_v_b_5_58483 = net_58483;
  assign seg_14_18_sp4_v_b_10_54660 = net_54660;
  assign seg_14_18_sp4_v_b_12_54772 = net_54772;
  assign seg_14_18_sp4_v_b_20_54780 = seg_14_16_sp4_v_b_44_54780;
  assign seg_14_18_sp4_v_b_2_54652 = seg_13_17_sp4_r_v_b_15_54652;
  assign seg_14_19_lutff_3_out_54997 = net_54997;
  assign seg_14_19_sp12_v_b_0_57482 = seg_14_13_sp12_v_b_12_57482;
  assign seg_14_19_sp12_v_b_10_58096 = seg_14_15_sp12_v_b_18_58096;
  assign seg_14_19_sp12_v_b_3_57605 = seg_14_14_sp12_v_b_12_57605;
  assign seg_14_19_sp4_v_b_22_54905 = net_54905;
  assign seg_14_1_neigh_op_lft_3_48911 = seg_13_1_lutff_3_out_48911;
  assign seg_14_1_neigh_op_tnl_0_49036 = seg_13_2_lutff_0_out_49036;
  assign seg_14_1_sp4_h_r_44_45228 = net_45228;
  assign seg_14_2_lutff_0_out_52867 = net_52867;
  assign seg_14_2_lutff_2_out_52869 = net_52869;
  assign seg_14_2_lutff_6_out_52873 = net_52873;
  assign seg_14_2_sp4_r_v_b_39_56883 = net_56883;
  assign seg_14_2_sp4_v_t_46_53183 = seg_13_4_sp4_r_v_b_35_53183;
  assign seg_14_3_lutff_6_out_53032 = net_53032;
  assign seg_14_3_lutff_7_out_53033 = net_53033;
  assign seg_14_3_sp4_h_l_41_41674 = seg_12_3_sp4_h_r_28_41674;
  assign seg_14_4_lutff_0_out_53149 = net_53149;
  assign seg_14_4_lutff_2_out_53151 = net_53151;
  assign seg_14_4_lutff_3_out_53152 = net_53152;
  assign seg_14_4_lutff_5_out_53154 = net_53154;
  assign seg_14_4_neigh_op_bnl_1_49196 = seg_13_3_lutff_1_out_49196;
  assign seg_14_4_neigh_op_bot_6_53032 = seg_14_3_lutff_6_out_53032;
  assign seg_14_4_neigh_op_bot_7_53033 = seg_14_3_lutff_7_out_53033;
  assign seg_14_4_neigh_op_lft_0_49318 = seg_13_4_lutff_0_out_49318;
  assign seg_14_4_sp4_h_r_20_53295 = net_53295;
  assign seg_14_4_sp4_h_r_30_49461 = net_49461;
  assign seg_14_4_sp4_h_r_36_45623 = net_45623;
  assign seg_14_4_sp4_r_v_b_15_56883 = seg_14_2_sp4_r_v_b_39_56883;
  assign seg_14_4_sp4_r_v_b_21_56889 = net_56889;
  assign seg_14_4_sp4_r_v_b_25_57003 = net_57003;
  assign seg_14_4_sp4_r_v_b_45_57135 = net_57135;
  assign seg_14_4_sp4_v_b_36_53296 = net_53296;
  assign seg_14_5_lutff_1_out_53273 = net_53273;
  assign seg_14_5_lutff_2_out_53274 = net_53274;
  assign seg_14_5_lutff_3_out_53275 = net_53275;
  assign seg_14_5_lutff_4_out_53276 = net_53276;
  assign seg_14_5_lutff_5_out_53277 = net_53277;
  assign seg_14_5_lutff_6_out_53278 = net_53278;
  assign seg_14_5_lutff_7_out_53279 = net_53279;
  assign seg_14_5_neigh_op_bnl_3_49321 = seg_13_4_lutff_3_out_49321;
  assign seg_14_5_neigh_op_bnl_4_49322 = seg_13_4_lutff_4_out_49322;
  assign seg_14_5_neigh_op_bot_0_53149 = seg_14_4_lutff_0_out_53149;
  assign seg_14_5_neigh_op_bot_3_53152 = seg_14_4_lutff_3_out_53152;
  assign seg_14_5_neigh_op_bot_5_53154 = seg_14_4_lutff_5_out_53154;
  assign seg_14_5_sp4_h_r_41_45751 = seg_11_5_sp4_h_r_4_45751;
  assign seg_14_5_sp4_r_v_b_17_57008 = net_57008;
  assign seg_14_5_sp4_v_b_11_53060 = seg_13_3_sp4_r_v_b_35_53060;
  assign seg_14_5_sp4_v_b_2_53053 = seg_13_4_sp4_r_v_b_15_53053;
  assign seg_14_6_lutff_0_out_53395 = net_53395;
  assign seg_14_6_lutff_3_out_53398 = net_53398;
  assign seg_14_6_lutff_5_out_53400 = net_53400;
  assign seg_14_6_lutff_7_out_53402 = net_53402;
  assign seg_14_6_neigh_op_bnl_0_49441 = seg_13_5_lutff_0_out_49441;
  assign seg_14_6_neigh_op_bot_3_53275 = seg_14_5_lutff_3_out_53275;
  assign seg_14_6_neigh_op_bot_7_53279 = seg_14_5_lutff_7_out_53279;
  assign seg_14_6_neigh_op_rgt_0_57225 = seg_15_6_lutff_0_out_57225;
  assign seg_14_6_neigh_op_rgt_4_57229 = seg_15_6_lutff_4_out_57229;
  assign seg_14_6_sp12_h_r_0_57356 = net_57356;
  assign seg_14_6_sp4_h_l_39_42041 = seg_10_6_sp4_h_r_2_42041;
  assign seg_14_6_sp4_h_l_42_42046 = seg_11_6_sp4_h_r_18_42046;
  assign seg_14_6_sp4_h_l_44_42048 = seg_13_6_sp4_h_r_44_42048;
  assign seg_14_6_sp4_h_r_0_57360 = seg_16_6_sp4_h_r_24_57360;
  assign seg_14_6_sp4_h_r_2_57364 = net_57364;
  assign seg_14_6_sp4_h_r_44_45879 = net_45879;
  assign seg_14_6_sp4_h_r_4_57366 = seg_16_6_sp4_h_r_28_57366;
  assign seg_14_6_sp4_h_r_8_57370 = net_57370;
  assign seg_14_6_sp4_r_v_b_1_57003 = seg_14_4_sp4_r_v_b_25_57003;
  assign seg_14_6_sp4_r_v_b_21_57135 = seg_14_4_sp4_r_v_b_45_57135;
  assign seg_14_6_sp4_v_b_12_53296 = seg_14_4_sp4_v_b_36_53296;
  assign seg_14_6_sp4_v_b_7_53179 = seg_13_6_sp4_r_v_b_7_53179;
  assign seg_14_7_lutff_1_out_53519 = net_53519;
  assign seg_14_7_lutff_5_out_53523 = net_53523;
  assign seg_14_7_lutff_6_out_53524 = net_53524;
  assign seg_14_7_lutff_7_out_53525 = net_53525;
  assign seg_14_7_neigh_op_bot_5_53400 = seg_14_6_lutff_5_out_53400;
  assign seg_14_7_neigh_op_rgt_2_57350 = seg_15_7_lutff_2_out_57350;
  assign seg_14_7_neigh_op_rgt_3_57351 = seg_15_7_lutff_3_out_57351;
  assign seg_14_7_sp4_h_l_37_42160 = seg_12_7_sp4_h_r_24_42160;
  assign seg_14_7_sp4_h_r_11_57486 = seg_17_7_sp4_h_r_46_57486;
  assign seg_14_7_sp4_h_r_12_53654 = net_53654;
  assign seg_14_7_sp4_h_r_28_49828 = net_49828;
  assign seg_14_7_sp4_h_r_38_45996 = net_45996;
  assign seg_14_7_sp4_v_b_1_53296 = seg_14_4_sp4_v_b_36_53296;
  assign seg_14_7_sp4_v_b_44_53673 = net_53673;
  assign seg_14_7_sp4_v_b_4_53301 = seg_13_4_sp4_r_v_b_41_53301;
  assign seg_14_8_lutff_5_out_53646 = net_53646;
  assign seg_14_8_neigh_op_bnl_0_49687 = seg_13_7_lutff_0_out_49687;
  assign seg_14_8_neigh_op_bnr_4_57352 = seg_15_7_lutff_4_out_57352;
  assign seg_14_8_neigh_op_bot_1_53519 = seg_14_7_lutff_1_out_53519;
  assign seg_14_8_neigh_op_bot_5_53523 = seg_14_7_lutff_5_out_53523;
  assign seg_14_8_neigh_op_top_0_53764 = seg_14_9_lutff_0_out_53764;
  assign seg_14_8_sp4_h_l_44_42294 = seg_11_8_sp4_h_r_20_42294;
  assign seg_14_8_sp4_h_r_0_57606 = net_57606;
  assign seg_14_8_sp4_h_r_11_57609 = seg_15_8_sp4_h_r_22_57609;
  assign seg_14_8_sp4_h_r_12_53777 = net_53777;
  assign seg_14_8_sp4_h_r_1_57607 = seg_17_8_sp4_h_r_36_57607;
  assign seg_14_8_sp4_h_r_22_53779 = net_53779;
  assign seg_14_8_sp4_h_r_2_57610 = net_57610;
  assign seg_14_8_sp4_h_r_38_46119 = net_46119;
  assign seg_14_8_sp4_h_r_40_46121 = net_46121;
  assign seg_14_8_sp4_h_r_46_46117 = net_46117;
  assign seg_14_8_sp4_h_r_5_57613 = seg_15_8_sp4_h_r_16_57613;
  assign seg_14_8_sp4_h_r_9_57617 = seg_17_8_sp4_h_r_44_57617;
  assign seg_14_8_sp4_r_v_b_39_57621 = net_57621;
  assign seg_14_8_sp4_r_v_b_47_57629 = net_57629;
  assign seg_14_8_sp4_v_b_20_53550 = net_53550;
  assign seg_14_8_sp4_v_b_22_53552 = net_53552;
  assign seg_14_8_sp4_v_b_32_53674 = seg_14_10_sp4_v_b_8_53674;
  assign seg_14_8_sp4_v_b_36_53788 = net_53788;
  assign seg_14_8_sp4_v_b_46_53798 = net_53798;
  assign seg_14_9_lutff_0_out_53764 = net_53764;
  assign seg_14_9_lutff_1_out_53765 = net_53765;
  assign seg_14_9_neigh_op_bnr_2_57473 = seg_15_8_lutff_2_out_57473;
  assign seg_14_9_neigh_op_bnr_4_57475 = seg_15_8_lutff_4_out_57475;
  assign seg_14_9_sp4_h_l_41_42412 = seg_12_9_sp4_h_r_28_42412;
  assign seg_14_9_sp4_h_l_45_42416 = seg_12_9_sp4_h_r_32_42416;
  assign seg_14_9_sp4_h_r_0_57729 = seg_16_9_sp4_h_r_24_57729;
  assign seg_14_9_sp4_h_r_10_57731 = seg_16_9_sp4_h_r_34_57731;
  assign seg_14_9_sp4_r_v_b_45_57750 = net_57750;
  assign seg_14_9_sp4_v_b_11_53552 = seg_14_8_sp4_v_b_22_53552;
  assign seg_14_9_sp4_v_b_17_53670 = seg_13_7_sp4_r_v_b_41_53670;
  assign seg_14_9_sp4_v_b_9_53550 = seg_14_8_sp4_v_b_20_53550;
  assign seg_15_0_span4_horz_r_0_60431 = seg_18_0_span4_horz_r_12_60431;
  assign seg_15_0_span4_vert_24_56738 = net_56738;
  assign seg_15_10_lutff_1_out_57718 = net_57718;
  assign seg_15_10_lutff_2_out_57719 = net_57719;
  assign seg_15_10_lutff_3_out_57720 = net_57720;
  assign seg_15_10_lutff_6_out_57723 = net_57723;
  assign seg_15_10_neigh_op_top_0_57840 = seg_15_11_lutff_0_out_57840;
  assign seg_15_10_sp4_h_r_0_61682 = seg_17_10_sp4_h_r_24_61682;
  assign seg_15_10_sp4_h_r_2_61686 = seg_17_10_sp4_h_r_26_61686;
  assign seg_15_10_sp4_h_r_30_54030 = net_54030;
  assign seg_15_10_sp4_v_b_8_57504 = seg_15_8_sp4_v_b_32_57504;
  assign seg_15_10_sp4_v_t_39_57990 = seg_15_12_sp4_v_b_26_57990;
  assign seg_15_11_lutff_0_out_57840 = net_57840;
  assign seg_15_11_lutff_1_out_57841 = net_57841;
  assign seg_15_11_lutff_2_out_57842 = net_57842;
  assign seg_15_11_lutff_3_out_57843 = net_57843;
  assign seg_15_11_lutff_4_out_57844 = net_57844;
  assign seg_15_11_lutff_7_out_57847 = net_57847;
  assign seg_15_11_neigh_op_bot_1_57718 = seg_15_10_lutff_1_out_57718;
  assign seg_15_11_neigh_op_bot_2_57719 = seg_15_10_lutff_2_out_57719;
  assign seg_15_11_neigh_op_bot_3_57720 = seg_15_10_lutff_3_out_57720;
  assign seg_15_11_neigh_op_bot_6_57723 = seg_15_10_lutff_6_out_57723;
  assign seg_15_11_neigh_op_rgt_6_61676 = seg_16_11_lutff_6_out_61676;
  assign seg_15_11_neigh_op_rgt_7_61677 = seg_16_11_lutff_7_out_61677;
  assign seg_15_11_sp4_h_r_0_61805 = net_61805;
  assign seg_15_11_sp4_h_r_16_57982 = net_57982;
  assign seg_15_11_sp4_h_r_22_57978 = net_57978;
  assign seg_15_11_sp4_h_r_28_54151 = net_54151;
  assign seg_15_11_sp4_h_r_42_50323 = net_50323;
  assign seg_15_11_sp4_h_r_5_61812 = seg_18_11_sp4_h_r_40_61812;
  assign seg_15_11_sp4_r_v_b_33_61702 = net_61702;
  assign seg_15_11_sp4_r_v_b_45_61826 = net_61826;
  assign seg_15_11_sp4_r_v_b_5_61452 = seg_16_8_sp4_v_b_40_61452;
  assign seg_15_11_sp4_v_b_0_57619 = seg_14_10_sp4_r_v_b_13_57619;
  assign seg_15_11_sp4_v_b_10_57629 = seg_14_8_sp4_r_v_b_47_57629;
  assign seg_15_11_sp4_v_b_12_57741 = net_57741;
  assign seg_15_11_sp4_v_b_2_57621 = seg_14_8_sp4_r_v_b_39_57621;
  assign seg_15_11_sp4_v_b_44_57995 = net_57995;
  assign seg_15_11_sp4_v_t_41_58115 = seg_15_13_sp4_v_b_28_58115;
  assign seg_15_12_lutff_1_out_57964 = net_57964;
  assign seg_15_12_lutff_2_out_57965 = net_57965;
  assign seg_15_12_lutff_3_out_57966 = net_57966;
  assign seg_15_12_lutff_4_out_57967 = net_57967;
  assign seg_15_12_lutff_6_out_57969 = net_57969;
  assign seg_15_12_lutff_7_out_57970 = net_57970;
  assign seg_15_12_neigh_op_bot_7_57847 = seg_15_11_lutff_7_out_57847;
  assign seg_15_12_neigh_op_top_7_58093 = seg_15_13_lutff_7_out_58093;
  assign seg_15_12_sp4_h_r_9_61939 = seg_16_12_sp4_h_r_20_61939;
  assign seg_15_12_sp4_r_v_b_33_61825 = net_61825;
  assign seg_15_12_sp4_r_v_b_47_61951 = seg_15_14_sp4_r_v_b_23_61951;
  assign seg_15_12_sp4_v_b_10_57752 = seg_14_11_sp4_r_v_b_23_57752;
  assign seg_15_12_sp4_v_b_11_57751 = seg_14_10_sp4_r_v_b_35_57751;
  assign seg_15_12_sp4_v_b_1_57741 = seg_15_11_sp4_v_b_12_57741;
  assign seg_15_12_sp4_v_b_25_57987 = seg_14_14_sp4_r_v_b_1_57987;
  assign seg_15_12_sp4_v_b_26_57990 = net_57990;
  assign seg_15_12_sp4_v_b_2_57744 = seg_14_11_sp4_r_v_b_15_57744;
  assign seg_15_12_sp4_v_b_34_57998 = seg_15_14_sp4_v_b_10_57998;
  assign seg_15_12_sp4_v_b_36_58110 = seg_15_14_sp4_v_b_12_58110;
  assign seg_15_12_sp4_v_b_3_57743 = seg_14_10_sp4_r_v_b_27_57743;
  assign seg_15_12_sp4_v_b_4_57746 = seg_14_11_sp4_r_v_b_17_57746;
  assign seg_15_12_sp4_v_b_5_57745 = seg_14_10_sp4_r_v_b_29_57745;
  assign seg_15_12_sp4_v_b_7_57747 = seg_14_10_sp4_r_v_b_31_57747;
  assign seg_15_12_sp4_v_b_8_57750 = seg_14_9_sp4_r_v_b_45_57750;
  assign seg_15_12_sp4_v_t_36_58233 = seg_15_15_sp4_v_b_12_58233;
  assign seg_15_13_lutff_1_out_58087 = net_58087;
  assign seg_15_13_lutff_2_out_58088 = net_58088;
  assign seg_15_13_lutff_3_out_58089 = net_58089;
  assign seg_15_13_lutff_5_out_58091 = net_58091;
  assign seg_15_13_lutff_7_out_58093 = net_58093;
  assign seg_15_13_neigh_op_rgt_1_61917 = seg_16_13_lutff_1_out_61917;
  assign seg_15_13_neigh_op_rgt_2_61918 = seg_16_13_lutff_2_out_61918;
  assign seg_15_13_neigh_op_rgt_3_61919 = seg_16_13_lutff_3_out_61919;
  assign seg_15_13_neigh_op_rgt_4_61920 = seg_16_13_lutff_4_out_61920;
  assign seg_15_13_neigh_op_rgt_5_61921 = seg_16_13_lutff_5_out_61921;
  assign seg_15_13_neigh_op_rgt_6_61922 = seg_16_13_lutff_6_out_61922;
  assign seg_15_13_neigh_op_top_5_58214 = seg_15_14_lutff_5_out_58214;
  assign seg_15_13_sp4_h_r_40_50567 = net_50567;
  assign seg_15_13_sp4_v_b_28_58115 = net_58115;
  assign seg_15_13_sp4_v_t_38_58358 = seg_14_17_sp4_r_v_b_3_58358;
  assign seg_15_14_lutff_1_out_58210 = net_58210;
  assign seg_15_14_lutff_4_out_58213 = net_58213;
  assign seg_15_14_lutff_5_out_58214 = net_58214;
  assign seg_15_14_neigh_op_bnl_0_54256 = seg_14_13_lutff_0_out_54256;
  assign seg_15_14_neigh_op_bot_1_58087 = seg_15_13_lutff_1_out_58087;
  assign seg_15_14_neigh_op_bot_2_58088 = seg_15_13_lutff_2_out_58088;
  assign seg_15_14_neigh_op_bot_3_58089 = seg_15_13_lutff_3_out_58089;
  assign seg_15_14_neigh_op_bot_5_58091 = seg_15_13_lutff_5_out_58091;
  assign seg_15_14_neigh_op_tnr_5_62167 = seg_16_15_lutff_5_out_62167;
  assign seg_15_14_neigh_op_top_4_58336 = seg_15_15_lutff_4_out_58336;
  assign seg_15_14_sp4_h_r_0_62174 = net_62174;
  assign seg_15_14_sp4_h_r_20_58355 = net_58355;
  assign seg_15_14_sp4_h_r_24_54514 = net_54514;
  assign seg_15_14_sp4_h_r_28_54520 = net_54520;
  assign seg_15_14_sp4_h_r_34_54516 = net_54516;
  assign seg_15_14_sp4_h_r_46_50686 = net_50686;
  assign seg_15_14_sp4_h_r_4_62180 = net_62180;
  assign seg_15_14_sp4_r_v_b_23_61951 = net_61951;
  assign seg_15_14_sp4_r_v_b_47_62197 = net_62197;
  assign seg_15_14_sp4_r_v_b_7_61823 = net_61823;
  assign seg_15_14_sp4_r_v_b_9_61825 = seg_15_12_sp4_r_v_b_33_61825;
  assign seg_15_14_sp4_v_b_10_57998 = net_57998;
  assign seg_15_14_sp4_v_b_12_58110 = net_58110;
  assign seg_15_14_sp4_v_b_8_57996 = seg_14_13_sp4_r_v_b_21_57996;
  assign seg_15_14_sp4_v_b_9_57995 = seg_15_11_sp4_v_b_44_57995;
  assign seg_15_14_sp4_v_t_43_58486 = seg_14_17_sp4_r_v_b_19_58486;
  assign seg_15_15_lutff_1_out_58333 = net_58333;
  assign seg_15_15_lutff_2_out_58334 = net_58334;
  assign seg_15_15_lutff_3_out_58335 = net_58335;
  assign seg_15_15_lutff_4_out_58336 = net_58336;
  assign seg_15_15_neigh_op_bot_1_58210 = seg_15_14_lutff_1_out_58210;
  assign seg_15_15_neigh_op_rgt_6_62168 = seg_16_15_lutff_6_out_62168;
  assign seg_15_15_sp4_h_l_44_46986 = seg_12_15_sp4_h_r_20_46986;
  assign seg_15_15_sp4_h_l_46_46978 = seg_12_15_sp4_h_r_22_46978;
  assign seg_15_15_sp4_r_v_b_15_62066 = net_62066;
  assign seg_15_15_sp4_r_v_b_17_62068 = net_62068;
  assign seg_15_15_sp4_r_v_b_9_61948 = net_61948;
  assign seg_15_15_sp4_v_b_12_58233 = net_58233;
  assign seg_15_15_sp4_v_b_32_58365 = net_58365;
  assign seg_15_15_sp4_v_b_45_58488 = seg_15_18_sp4_v_b_8_58488;
  assign seg_15_15_sp4_v_b_7_58116 = seg_14_13_sp4_r_v_b_31_58116;
  assign seg_15_16_lutff_1_out_58456 = net_58456;
  assign seg_15_16_lutff_2_out_58457 = net_58457;
  assign seg_15_16_lutff_4_out_58459 = net_58459;
  assign seg_15_16_lutff_5_out_58460 = net_58460;
  assign seg_15_16_lutff_7_out_58462 = net_58462;
  assign seg_15_16_neigh_op_rgt_0_62285 = seg_16_16_lutff_0_out_62285;
  assign seg_15_16_neigh_op_rgt_1_62286 = seg_16_16_lutff_1_out_62286;
  assign seg_15_16_neigh_op_rgt_6_62291 = seg_16_16_lutff_6_out_62291;
  assign seg_15_16_neigh_op_tnr_2_62410 = seg_16_17_lutff_2_out_62410;
  assign seg_15_16_sp4_v_b_11_58243 = seg_14_16_sp4_r_v_b_11_58243;
  assign seg_15_16_sp4_v_b_13_58357 = seg_14_14_sp4_r_v_b_37_58357;
  assign seg_15_16_sp4_v_b_17_58361 = seg_14_14_sp4_r_v_b_41_58361;
  assign seg_15_16_sp4_v_b_19_58363 = seg_14_14_sp4_r_v_b_43_58363;
  assign seg_15_16_sp4_v_b_23_58367 = seg_14_14_sp4_r_v_b_47_58367;
  assign seg_15_16_sp4_v_b_27_58481 = seg_14_18_sp4_r_v_b_3_58481;
  assign seg_15_16_sp4_v_b_29_58483 = seg_14_18_sp4_r_v_b_5_58483;
  assign seg_15_16_sp4_v_b_2_58236 = seg_14_13_sp4_r_v_b_39_58236;
  assign seg_15_16_sp4_v_b_35_58489 = seg_14_18_sp4_r_v_b_11_58489;
  assign seg_15_16_sp4_v_b_37_58603 = seg_14_18_sp4_r_v_b_13_58603;
  assign seg_15_16_sp4_v_b_38_58604 = net_58604;
  assign seg_15_16_sp4_v_b_44_58610 = net_58610;
  assign seg_15_16_sp4_v_b_9_58241 = seg_14_14_sp4_r_v_b_33_58241;
  assign seg_15_17_lutff_0_out_58578 = net_58578;
  assign seg_15_17_lutff_2_out_58580 = net_58580;
  assign seg_15_17_lutff_4_out_58582 = net_58582;
  assign seg_15_17_neigh_op_rgt_3_62411 = seg_16_17_lutff_3_out_62411;
  assign seg_15_17_neigh_op_tnl_1_54872 = seg_14_18_lutff_1_out_54872;
  assign seg_15_17_neigh_op_tnl_5_54876 = seg_14_18_lutff_5_out_54876;
  assign seg_15_17_neigh_op_tnl_7_54878 = seg_14_18_lutff_7_out_54878;
  assign seg_15_17_sp4_h_r_0_62543 = seg_17_17_sp4_h_r_24_62543;
  assign seg_15_17_sp4_h_r_16_58720 = seg_17_17_sp4_h_r_40_58720;
  assign seg_15_17_sp4_h_r_2_62547 = net_62547;
  assign seg_15_17_sp4_v_b_6_58363 = seg_14_14_sp4_r_v_b_43_58363;
  assign seg_15_17_sp4_v_b_8_58365 = seg_15_15_sp4_v_b_32_58365;
  assign seg_15_18_sp4_v_b_8_58488 = net_58488;
  assign seg_15_1_sp4_h_l_44_45228 = seg_14_1_sp4_h_r_44_45228;
  assign seg_15_2_sp4_h_l_47_45378 = seg_11_2_sp4_h_r_10_45378;
  assign seg_15_2_sp4_h_r_11_60701 = seg_16_2_sp4_h_r_22_60701;
  assign seg_15_2_sp4_h_r_39_49211 = seg_12_2_sp4_h_r_2_49211;
  assign seg_15_2_sp4_h_r_5_60705 = seg_18_2_sp4_h_r_40_60705;
  assign seg_15_2_sp4_v_b_28_56757 = net_56757;
  assign seg_15_3_lutff_2_out_56858 = net_56858;
  assign seg_15_3_neigh_op_top_2_56981 = seg_15_4_lutff_2_out_56981;
  assign seg_15_3_sp4_h_r_12_56992 = seg_17_3_sp4_h_r_36_56992;
  assign seg_15_3_sp4_h_r_40_49337 = net_49337;
  assign seg_15_3_sp4_v_b_0_56738 = seg_15_0_span4_vert_24_56738;
  assign seg_15_4_lutff_0_out_56979 = net_56979;
  assign seg_15_4_lutff_2_out_56981 = net_56981;
  assign seg_15_4_lutff_7_out_56986 = net_56986;
  assign seg_15_4_neigh_op_lft_2_53151 = seg_14_4_lutff_2_out_53151;
  assign seg_15_4_sp4_h_r_24_53284 = net_53284;
  assign seg_15_4_sp4_h_r_26_53288 = net_53288;
  assign seg_15_4_sp4_h_r_28_53290 = seg_13_4_sp4_h_r_4_53290;
  assign seg_15_4_sp4_h_r_32_53294 = seg_13_4_sp4_h_r_8_53294;
  assign seg_15_4_sp4_h_r_34_53286 = net_53286;
  assign seg_15_4_sp4_h_r_40_49460 = seg_13_4_sp4_h_r_16_49460;
  assign seg_15_4_sp4_h_r_6_60952 = net_60952;
  assign seg_15_4_sp4_r_v_b_29_60837 = net_60837;
  assign seg_15_4_sp4_r_v_b_39_60959 = net_60959;
  assign seg_15_4_sp4_r_v_b_41_60961 = net_60961;
  assign seg_15_4_sp4_v_b_36_57126 = seg_15_6_sp4_v_b_12_57126;
  assign seg_15_4_sp4_v_b_44_57134 = net_57134;
  assign seg_15_4_sp4_v_b_4_56757 = seg_15_2_sp4_v_b_28_56757;
  assign seg_15_4_sp4_v_t_37_57250 = seg_15_8_sp4_v_b_0_57250;
  assign seg_15_5_neigh_op_bnl_2_53151 = seg_14_4_lutff_2_out_53151;
  assign seg_15_5_sp12_v_b_4_60411 = net_60411;
  assign seg_15_5_sp4_h_l_41_45751 = seg_11_5_sp4_h_r_4_45751;
  assign seg_15_5_sp4_h_l_47_45747 = seg_11_5_sp4_h_r_10_45747;
  assign seg_15_5_sp4_h_r_24_53407 = net_53407;
  assign seg_15_5_sp4_h_r_26_53411 = net_53411;
  assign seg_15_5_sp4_h_r_30_53415 = net_53415;
  assign seg_15_5_sp4_r_v_b_13_60834 = net_60834;
  assign seg_15_5_sp4_r_v_b_21_60842 = net_60842;
  assign seg_15_5_sp4_r_v_b_23_60844 = net_60844;
  assign seg_15_5_sp4_r_v_b_29_60960 = net_60960;
  assign seg_15_5_sp4_r_v_b_33_60964 = net_60964;
  assign seg_15_5_sp4_v_b_16_57007 = net_57007;
  assign seg_15_5_sp4_v_b_18_57009 = net_57009;
  assign seg_15_5_sp4_v_b_34_57137 = net_57137;
  assign seg_15_5_sp4_v_b_8_56889 = seg_14_4_sp4_r_v_b_21_56889;
  assign seg_15_6_lutff_0_out_57225 = net_57225;
  assign seg_15_6_lutff_4_out_57229 = net_57229;
  assign seg_15_6_lutff_7_out_57232 = net_57232;
  assign seg_15_6_neigh_op_bnl_4_53276 = seg_14_5_lutff_4_out_53276;
  assign seg_15_6_neigh_op_bnl_5_53277 = seg_14_5_lutff_5_out_53277;
  assign seg_15_6_neigh_op_lft_3_53398 = seg_14_6_lutff_3_out_53398;
  assign seg_15_6_neigh_op_lft_7_53402 = seg_14_6_lutff_7_out_53402;
  assign seg_15_6_sp4_h_l_39_45872 = seg_11_6_sp4_h_r_2_45872;
  assign seg_15_6_sp4_h_l_43_45876 = seg_13_6_sp4_h_r_30_45876;
  assign seg_15_6_sp4_h_r_26_53534 = seg_13_6_sp4_h_r_2_53534;
  assign seg_15_6_sp4_h_r_2_61194 = net_61194;
  assign seg_15_6_sp4_h_r_32_53540 = seg_13_6_sp4_h_r_8_53540;
  assign seg_15_6_sp4_h_r_38_49704 = net_49704;
  assign seg_15_6_sp4_h_r_42_49708 = net_49708;
  assign seg_15_6_sp4_h_r_44_49710 = seg_13_6_sp4_h_r_20_49710;
  assign seg_15_6_sp4_h_r_9_61201 = seg_16_6_sp4_h_r_20_61201;
  assign seg_15_6_sp4_v_b_12_57126 = net_57126;
  assign seg_15_6_sp4_v_b_4_57008 = seg_14_5_sp4_r_v_b_17_57008;
  assign seg_15_6_sp4_v_b_5_57007 = seg_15_5_sp4_v_b_16_57007;
  assign seg_15_6_sp4_v_b_7_57009 = seg_15_5_sp4_v_b_18_57009;
  assign seg_15_7_lutff_2_out_57350 = net_57350;
  assign seg_15_7_lutff_3_out_57351 = net_57351;
  assign seg_15_7_lutff_4_out_57352 = net_57352;
  assign seg_15_7_lutff_6_out_57354 = net_57354;
  assign seg_15_7_neigh_op_bot_7_57232 = seg_15_6_lutff_7_out_57232;
  assign seg_15_7_sp12_v_b_0_60411 = seg_15_5_sp12_v_b_4_60411;
  assign seg_15_7_sp4_h_l_37_45991 = seg_11_7_sp4_h_r_0_45991;
  assign seg_15_7_sp4_h_l_47_45993 = seg_11_7_sp4_h_r_10_45993;
  assign seg_15_7_sp4_h_r_5_61320 = seg_18_7_sp4_h_r_40_61320;
  assign seg_15_7_sp4_h_r_7_61322 = seg_18_7_sp4_h_r_42_61322;
  assign seg_15_7_sp4_h_r_9_61324 = seg_16_7_sp4_h_r_20_61324;
  assign seg_15_7_sp4_v_b_10_57137 = seg_15_5_sp4_v_b_34_57137;
  assign seg_15_7_sp4_v_b_9_57134 = seg_15_4_sp4_v_b_44_57134;
  assign seg_15_7_sp4_v_t_36_57618 = seg_15_8_sp4_v_b_36_57618;
  assign seg_15_8_lutff_2_out_57473 = net_57473;
  assign seg_15_8_lutff_3_out_57474 = net_57474;
  assign seg_15_8_lutff_4_out_57475 = net_57475;
  assign seg_15_8_neigh_op_lft_5_53646 = seg_14_8_lutff_5_out_53646;
  assign seg_15_8_neigh_op_rgt_0_61301 = seg_16_8_lutff_0_out_61301;
  assign seg_15_8_sp4_h_l_45_46124 = seg_13_8_sp4_h_r_32_46124;
  assign seg_15_8_sp4_h_r_10_61438 = seg_17_8_sp4_h_r_34_61438;
  assign seg_15_8_sp4_h_r_11_61439 = seg_18_8_sp4_h_r_46_61439;
  assign seg_15_8_sp4_h_r_16_57613 = net_57613;
  assign seg_15_8_sp4_h_r_22_57609 = net_57609;
  assign seg_15_8_sp4_h_r_24_53776 = net_53776;
  assign seg_15_8_sp4_h_r_34_53778 = net_53778;
  assign seg_15_8_sp4_h_r_40_49952 = net_49952;
  assign seg_15_8_sp4_h_r_5_61443 = seg_18_8_sp4_h_r_40_61443;
  assign seg_15_8_sp4_r_v_b_23_61213 = net_61213;
  assign seg_15_8_sp4_r_v_b_35_61335 = net_61335;
  assign seg_15_8_sp4_r_v_b_3_61081 = net_61081;
  assign seg_15_8_sp4_v_b_0_57250 = net_57250;
  assign seg_15_8_sp4_v_b_32_57504 = net_57504;
  assign seg_15_8_sp4_v_b_36_57618 = net_57618;
  assign seg_15_9_neigh_op_bot_2_57473 = seg_15_8_lutff_2_out_57473;
  assign seg_15_9_neigh_op_bot_3_57474 = seg_15_8_lutff_3_out_57474;
  assign seg_15_9_neigh_op_bot_4_57475 = seg_15_8_lutff_4_out_57475;
  assign seg_15_9_neigh_op_rgt_4_61428 = seg_16_9_lutff_4_out_61428;
  assign seg_15_9_neigh_op_rgt_7_61431 = seg_16_9_lutff_7_out_61431;
  assign seg_15_9_sp4_h_r_28_53905 = net_53905;
  assign seg_15_9_sp4_h_r_32_53909 = net_53909;
  assign seg_15_9_sp4_r_v_b_37_61572 = net_61572;
  assign seg_15_9_sp4_r_v_b_39_61574 = net_61574;
  assign seg_15_9_sp4_r_v_b_3_61204 = net_61204;
  assign seg_15_9_sp4_r_v_b_41_61576 = net_61576;
  assign seg_16_0_span4_horz_r_0_64262 = seg_19_0_span4_horz_r_12_64262;
  assign seg_16_10_lutff_1_out_61548 = net_61548;
  assign seg_16_10_neigh_op_rgt_1_65379 = seg_17_10_lutff_1_out_65379;
  assign seg_16_10_neigh_op_tnl_3_57843 = seg_15_11_lutff_3_out_57843;
  assign seg_16_10_sp4_r_v_b_17_65284 = net_65284;
  assign seg_16_10_sp4_r_v_b_21_65288 = net_65288;
  assign seg_16_10_sp4_r_v_b_23_65290 = net_65290;
  assign seg_16_10_sp4_r_v_b_29_65406 = net_65406;
  assign seg_16_10_sp4_r_v_b_31_65408 = net_65408;
  assign seg_16_10_sp4_r_v_b_33_65410 = net_65410;
  assign seg_16_10_sp4_r_v_b_39_65528 = net_65528;
  assign seg_16_10_sp4_r_v_b_41_65530 = net_65530;
  assign seg_16_10_sp4_r_v_b_43_65532 = net_65532;
  assign seg_16_10_sp4_v_b_10_61336 = seg_16_8_sp4_v_b_34_61336;
  assign seg_16_10_sp4_v_b_11_61335 = seg_15_8_sp4_r_v_b_35_61335;
  assign seg_16_10_sp4_v_t_42_61823 = seg_15_14_sp4_r_v_b_7_61823;
  assign seg_16_11_lutff_1_out_61671 = net_61671;
  assign seg_16_11_lutff_3_out_61673 = net_61673;
  assign seg_16_11_lutff_5_out_61675 = net_61675;
  assign seg_16_11_lutff_6_out_61676 = net_61676;
  assign seg_16_11_lutff_7_out_61677 = net_61677;
  assign seg_16_11_neigh_op_bnr_5_65383 = seg_17_10_lutff_5_out_65383;
  assign seg_16_11_neigh_op_bot_1_61548 = seg_16_10_lutff_1_out_61548;
  assign seg_16_11_neigh_op_rgt_1_65502 = seg_17_11_lutff_1_out_65502;
  assign seg_16_11_neigh_op_rgt_2_65503 = seg_17_11_lutff_2_out_65503;
  assign seg_16_11_neigh_op_rgt_3_65504 = seg_17_11_lutff_3_out_65504;
  assign seg_16_11_neigh_op_rgt_4_65505 = seg_17_11_lutff_4_out_65505;
  assign seg_16_11_neigh_op_tnl_6_57969 = seg_15_12_lutff_6_out_57969;
  assign seg_16_11_sp12_v_b_18_65265 = net_65265;
  assign seg_16_11_sp12_v_b_22_65511 = net_65511;
  assign seg_16_11_sp4_h_l_37_50314 = seg_14_11_sp4_h_r_24_50314;
  assign seg_16_11_sp4_h_l_41_50320 = seg_12_11_sp4_h_r_4_50320;
  assign seg_16_11_sp4_h_r_0_65636 = seg_18_11_sp4_h_r_24_65636;
  assign seg_16_11_sp4_h_r_24_57975 = net_57975;
  assign seg_16_11_sp4_h_r_36_54146 = net_54146;
  assign seg_16_11_sp4_h_r_8_65646 = net_65646;
  assign seg_16_11_sp4_r_v_b_21_65411 = net_65411;
  assign seg_16_11_sp4_v_b_10_61459 = seg_16_9_sp4_v_b_34_61459;
  assign seg_16_11_sp4_v_b_12_61571 = net_61571;
  assign seg_16_11_sp4_v_b_14_61573 = net_61573;
  assign seg_16_12_sp4_h_l_43_50445 = seg_12_12_sp4_h_r_6_50445;
  assign seg_16_12_sp4_h_r_12_61929 = net_61929;
  assign seg_16_12_sp4_h_r_20_61939 = net_61939;
  assign seg_16_12_sp4_h_r_30_58106 = net_58106;
  assign seg_16_12_sp4_v_b_0_61572 = seg_15_9_sp4_r_v_b_37_61572;
  assign seg_16_12_sp4_v_b_4_61576 = seg_15_9_sp4_r_v_b_41_61576;
  assign seg_16_12_sp4_v_b_6_61578 = net_61578;
  assign seg_16_12_sp4_v_b_7_61577 = seg_16_9_sp4_v_b_42_61577;
  assign seg_16_13_lutff_1_out_61917 = net_61917;
  assign seg_16_13_lutff_2_out_61918 = net_61918;
  assign seg_16_13_lutff_3_out_61919 = net_61919;
  assign seg_16_13_lutff_4_out_61920 = net_61920;
  assign seg_16_13_lutff_5_out_61921 = net_61921;
  assign seg_16_13_lutff_6_out_61922 = net_61922;
  assign seg_16_13_neigh_op_bnl_2_57965 = seg_15_12_lutff_2_out_57965;
  assign seg_16_13_neigh_op_bnl_3_57966 = seg_15_12_lutff_3_out_57966;
  assign seg_16_13_neigh_op_bnl_4_57967 = seg_15_12_lutff_4_out_57967;
  assign seg_16_13_sp12_v_b_11_65020 = seg_16_18_sp12_v_b_0_65020;
  assign seg_16_13_sp4_h_l_40_50567 = seg_15_13_sp4_h_r_40_50567;
  assign seg_16_13_sp4_h_r_10_65884 = seg_18_13_sp4_h_r_34_65884;
  assign seg_16_13_sp4_h_r_12_62052 = seg_18_13_sp4_h_r_36_62052;
  assign seg_16_13_sp4_h_r_16_62058 = seg_18_13_sp4_h_r_40_62058;
  assign seg_16_13_sp4_h_r_20_62062 = seg_18_13_sp4_h_r_44_62062;
  assign seg_16_13_sp4_h_r_24_58221 = seg_14_13_sp4_h_r_0_58221;
  assign seg_16_13_sp4_h_r_34_58223 = seg_14_13_sp4_h_r_10_58223;
  assign seg_16_13_sp4_r_v_b_15_65651 = net_65651;
  assign seg_16_13_sp4_r_v_b_31_65777 = net_65777;
  assign seg_16_13_sp4_v_b_33_61948 = seg_15_15_sp4_r_v_b_9_61948;
  assign seg_16_13_sp4_v_b_39_62066 = seg_15_15_sp4_r_v_b_15_62066;
  assign seg_16_13_sp4_v_b_46_62073 = seg_16_15_sp4_v_b_22_62073;
  assign seg_16_13_sp4_v_b_9_61702 = seg_15_11_sp4_r_v_b_33_61702;
  assign seg_16_13_sp4_v_t_43_62193 = seg_16_17_sp4_v_b_6_62193;
  assign seg_16_13_sp4_v_t_47_62197 = seg_15_14_sp4_r_v_b_47_62197;
  assign seg_16_14_lutff_1_out_62040 = net_62040;
  assign seg_16_14_lutff_2_out_62041 = net_62041;
  assign seg_16_14_lutff_3_out_62042 = net_62042;
  assign seg_16_14_lutff_4_out_62043 = net_62043;
  assign seg_16_14_lutff_5_out_62044 = net_62044;
  assign seg_16_14_lutff_6_out_62045 = net_62045;
  assign seg_16_14_lutff_7_out_62046 = net_62046;
  assign seg_16_14_neigh_op_rgt_5_65875 = seg_17_14_lutff_5_out_65875;
  assign seg_16_14_neigh_op_tnl_3_58335 = seg_15_15_lutff_3_out_58335;
  assign seg_16_14_neigh_op_tnr_0_65993 = seg_17_15_lutff_0_out_65993;
  assign seg_16_14_neigh_op_tnr_2_65995 = seg_17_15_lutff_2_out_65995;
  assign seg_16_14_neigh_op_tnr_3_65996 = seg_17_15_lutff_3_out_65996;
  assign seg_16_14_neigh_op_tnr_7_66000 = seg_17_15_lutff_7_out_66000;
  assign seg_16_14_neigh_op_top_1_62163 = seg_16_15_lutff_1_out_62163;
  assign seg_16_14_neigh_op_top_2_62164 = seg_16_15_lutff_2_out_62164;
  assign seg_16_14_neigh_op_top_7_62169 = seg_16_15_lutff_7_out_62169;
  assign seg_16_14_sp4_h_l_42_50692 = seg_13_14_sp4_h_r_18_50692;
  assign seg_16_14_sp4_h_l_43_50691 = seg_14_14_sp4_h_r_30_50691;
  assign seg_16_14_sp4_h_l_46_50686 = seg_15_14_sp4_h_r_46_50686;
  assign seg_16_14_sp4_h_r_12_62175 = seg_18_14_sp4_h_r_36_62175;
  assign seg_16_14_sp4_h_r_13_62174 = seg_15_14_sp4_h_r_0_62174;
  assign seg_16_14_sp4_h_r_14_62179 = seg_18_14_sp4_h_r_38_62179;
  assign seg_16_14_sp4_h_r_16_62181 = seg_18_14_sp4_h_r_40_62181;
  assign seg_16_14_sp4_h_r_6_66013 = seg_18_14_sp4_h_r_30_66013;
  assign seg_16_14_sp4_h_r_8_66015 = seg_18_14_sp4_h_r_32_66015;
  assign seg_16_14_sp4_v_b_8_61826 = seg_15_11_sp4_r_v_b_45_61826;
  assign seg_16_15_lutff_0_out_62162 = net_62162;
  assign seg_16_15_lutff_1_out_62163 = net_62163;
  assign seg_16_15_lutff_2_out_62164 = net_62164;
  assign seg_16_15_lutff_4_out_62166 = net_62166;
  assign seg_16_15_lutff_5_out_62167 = net_62167;
  assign seg_16_15_lutff_6_out_62168 = net_62168;
  assign seg_16_15_lutff_7_out_62169 = net_62169;
  assign seg_16_15_neigh_op_bnr_7_65877 = seg_17_14_lutff_7_out_65877;
  assign seg_16_15_neigh_op_rgt_1_65994 = seg_17_15_lutff_1_out_65994;
  assign seg_16_15_neigh_op_rgt_5_65998 = seg_17_15_lutff_5_out_65998;
  assign seg_16_15_neigh_op_rgt_6_65999 = seg_17_15_lutff_6_out_65999;
  assign seg_16_15_neigh_op_top_7_62292 = seg_16_16_lutff_7_out_62292;
  assign seg_16_15_sp4_h_l_37_50806 = seg_12_15_sp4_h_r_0_50806;
  assign seg_16_15_sp4_h_l_41_50812 = seg_12_15_sp4_h_r_4_50812;
  assign seg_16_15_sp4_h_r_10_66130 = net_66130;
  assign seg_16_15_sp4_h_r_12_62298 = net_62298;
  assign seg_16_15_sp4_h_r_24_58467 = net_58467;
  assign seg_16_15_sp4_r_v_b_11_65781 = net_65781;
  assign seg_16_15_sp4_v_b_22_62073 = net_62073;
  assign seg_16_15_sp4_v_b_24_62187 = seg_16_17_sp4_v_b_0_62187;
  assign seg_16_16_lutff_0_out_62285 = net_62285;
  assign seg_16_16_lutff_1_out_62286 = net_62286;
  assign seg_16_16_lutff_2_out_62287 = net_62287;
  assign seg_16_16_lutff_3_out_62288 = net_62288;
  assign seg_16_16_lutff_4_out_62289 = net_62289;
  assign seg_16_16_lutff_6_out_62291 = net_62291;
  assign seg_16_16_lutff_7_out_62292 = net_62292;
  assign seg_16_16_neigh_op_lft_2_58457 = seg_15_16_lutff_2_out_58457;
  assign seg_16_16_neigh_op_lft_4_58459 = seg_15_16_lutff_4_out_58459;
  assign seg_16_16_neigh_op_lft_5_58460 = seg_15_16_lutff_5_out_58460;
  assign seg_16_16_neigh_op_lft_7_58462 = seg_15_16_lutff_7_out_58462;
  assign seg_16_16_neigh_op_top_0_62408 = seg_16_17_lutff_0_out_62408;
  assign seg_16_16_sp4_h_l_37_50929 = seg_14_16_sp4_h_r_24_50929;
  assign seg_16_16_sp4_h_l_46_50932 = seg_13_16_sp4_h_r_22_50932;
  assign seg_16_16_sp4_h_r_10_66253 = seg_18_16_sp4_h_r_34_66253;
  assign seg_16_16_sp4_h_r_28_58596 = seg_14_16_sp4_h_r_4_58596;
  assign seg_16_16_sp4_h_r_32_58600 = net_58600;
  assign seg_16_16_sp4_h_r_34_58592 = net_58592;
  assign seg_16_16_sp4_h_r_38_54765 = seg_14_16_sp4_h_r_14_54765;
  assign seg_16_16_sp4_h_r_44_54771 = net_54771;
  assign seg_16_16_sp4_h_r_8_66261 = net_66261;
  assign seg_16_16_sp4_r_v_b_11_65904 = net_65904;
  assign seg_16_16_sp4_v_b_4_62068 = seg_15_15_sp4_r_v_b_17_62068;
  assign seg_16_16_sp4_v_t_36_62555 = seg_16_17_sp4_v_b_36_62555;
  assign seg_16_17_lutff_0_out_62408 = net_62408;
  assign seg_16_17_lutff_1_out_62409 = net_62409;
  assign seg_16_17_lutff_2_out_62410 = net_62410;
  assign seg_16_17_lutff_3_out_62411 = net_62411;
  assign seg_16_17_lutff_4_out_62412 = net_62412;
  assign seg_16_17_lutff_5_out_62413 = net_62413;
  assign seg_16_17_lutff_6_out_62414 = net_62414;
  assign seg_16_17_neigh_op_bnl_1_58456 = seg_15_16_lutff_1_out_58456;
  assign seg_16_17_neigh_op_lft_0_58578 = seg_15_17_lutff_0_out_58578;
  assign seg_16_17_neigh_op_lft_4_58582 = seg_15_17_lutff_4_out_58582;
  assign seg_16_17_neigh_op_tnr_6_66368 = seg_17_18_lutff_6_out_66368;
  assign seg_16_17_sp4_h_l_38_51057 = seg_13_17_sp4_h_r_14_51057;
  assign seg_16_17_sp4_h_r_14_62548 = net_62548;
  assign seg_16_17_sp4_h_r_24_58713 = seg_14_17_sp4_h_r_0_58713;
  assign seg_16_17_sp4_h_r_38_54888 = net_54888;
  assign seg_16_17_sp4_h_r_3_66379 = seg_17_17_sp4_h_r_14_66379;
  assign seg_16_17_sp4_r_v_b_13_66141 = net_66141;
  assign seg_16_17_sp4_r_v_b_3_66019 = net_66019;
  assign seg_16_17_sp4_r_v_b_43_66393 = net_66393;
  assign seg_16_17_sp4_r_v_b_9_66025 = net_66025;
  assign seg_16_17_sp4_v_b_0_62187 = net_62187;
  assign seg_16_17_sp4_v_b_36_62555 = net_62555;
  assign seg_16_17_sp4_v_b_6_62193 = net_62193;
  assign seg_16_18_sp12_v_b_0_65020 = net_65020;
  assign seg_16_1_sp4_h_l_46_49051 = seg_13_1_sp4_h_r_22_49051;
  assign seg_16_20_sp12_v_b_1_65265 = seg_16_11_sp12_v_b_18_65265;
  assign seg_16_22_sp12_v_b_1_65511 = seg_16_11_sp12_v_b_22_65511;
  assign seg_16_2_sp4_h_l_39_49211 = seg_12_2_sp4_h_r_2_49211;
  assign seg_16_2_sp4_h_r_0_64529 = seg_18_2_sp4_h_r_24_64529;
  assign seg_16_2_sp4_h_r_22_60701 = net_60701;
  assign seg_16_2_sp4_v_t_47_60844 = seg_15_5_sp4_r_v_b_23_60844;
  assign seg_16_3_lutff_2_out_60688 = net_60688;
  assign seg_16_3_sp12_v_b_4_64260 = net_64260;
  assign seg_16_3_sp4_h_r_36_53162 = net_53162;
  assign seg_16_3_sp4_h_r_4_64658 = net_64658;
  assign seg_16_3_sp4_h_r_6_64660 = net_64660;
  assign seg_16_3_sp4_r_v_b_23_64424 = net_64424;
  assign seg_16_3_sp4_r_v_b_37_64665 = net_64665;
  assign seg_16_3_sp4_v_b_20_60590 = net_60590;
  assign seg_16_3_sp4_v_b_36_60833 = net_60833;
  assign seg_16_3_sp4_v_b_38_60835 = net_60835;
  assign seg_16_4_neigh_op_bnl_2_56858 = seg_15_3_lutff_2_out_56858;
  assign seg_16_4_neigh_op_bnr_3_64520 = seg_17_3_lutff_3_out_64520;
  assign seg_16_4_neigh_op_bnr_4_64521 = seg_17_3_lutff_4_out_64521;
  assign seg_16_4_neigh_op_lft_7_56986 = seg_15_4_lutff_7_out_56986;
  assign seg_16_4_neigh_op_rgt_0_64640 = seg_17_4_lutff_0_out_64640;
  assign seg_16_4_neigh_op_rgt_1_64641 = seg_17_4_lutff_1_out_64641;
  assign seg_16_4_neigh_op_rgt_3_64643 = seg_17_4_lutff_3_out_64643;
  assign seg_16_4_neigh_op_rgt_4_64644 = seg_17_4_lutff_4_out_64644;
  assign seg_16_4_neigh_op_rgt_5_64645 = seg_17_4_lutff_5_out_64645;
  assign seg_16_4_neigh_op_rgt_6_64646 = seg_17_4_lutff_6_out_64646;
  assign seg_16_4_neigh_op_rgt_7_64647 = seg_17_4_lutff_7_out_64647;
  assign seg_16_4_neigh_op_tnr_0_64763 = seg_17_5_lutff_0_out_64763;
  assign seg_16_4_neigh_op_tnr_6_64769 = seg_17_5_lutff_6_out_64769;
  assign seg_16_4_neigh_op_top_4_60936 = seg_16_5_lutff_4_out_60936;
  assign seg_16_4_neigh_op_top_6_60938 = seg_16_5_lutff_6_out_60938;
  assign seg_16_4_neigh_op_top_7_60939 = seg_16_5_lutff_7_out_60939;
  assign seg_16_4_sp4_r_v_b_27_64666 = net_64666;
  assign seg_16_4_sp4_r_v_b_35_64674 = net_64674;
  assign seg_16_4_sp4_r_v_b_41_64792 = net_64792;
  assign seg_16_4_sp4_r_v_b_45_64796 = net_64796;
  assign seg_16_4_sp4_v_b_36_60956 = net_60956;
  assign seg_16_4_sp4_v_b_38_60958 = net_60958;
  assign seg_16_4_sp4_v_b_46_60966 = net_60966;
  assign seg_16_4_sp4_v_b_9_60590 = seg_16_3_sp4_v_b_20_60590;
  assign seg_16_4_sp4_v_t_38_61081 = seg_15_8_sp4_r_v_b_3_61081;
  assign seg_16_5_lutff_4_out_60936 = net_60936;
  assign seg_16_5_lutff_5_out_60937 = net_60937;
  assign seg_16_5_lutff_6_out_60938 = net_60938;
  assign seg_16_5_lutff_7_out_60939 = net_60939;
  assign seg_16_5_neigh_op_rgt_0_64763 = seg_17_5_lutff_0_out_64763;
  assign seg_16_5_neigh_op_rgt_1_64764 = seg_17_5_lutff_1_out_64764;
  assign seg_16_5_neigh_op_rgt_2_64765 = seg_17_5_lutff_2_out_64765;
  assign seg_16_5_neigh_op_rgt_3_64766 = seg_17_5_lutff_3_out_64766;
  assign seg_16_5_neigh_op_rgt_6_64769 = seg_17_5_lutff_6_out_64769;
  assign seg_16_5_neigh_op_rgt_7_64770 = seg_17_5_lutff_7_out_64770;
  assign seg_16_5_neigh_op_tnr_2_64888 = seg_17_6_lutff_2_out_64888;
  assign seg_16_5_neigh_op_tnr_6_64892 = seg_17_6_lutff_6_out_64892;
  assign seg_16_5_sp12_v_b_0_64260 = seg_16_3_sp12_v_b_4_64260;
  assign seg_16_5_sp4_h_l_37_49576 = seg_12_5_sp4_h_r_0_49576;
  assign seg_16_5_sp4_h_l_47_49578 = seg_12_5_sp4_h_r_10_49578;
  assign seg_16_5_sp4_r_v_b_39_64913 = net_64913;
  assign seg_16_5_sp4_v_b_32_60965 = net_60965;
  assign seg_16_5_sp4_v_b_34_60967 = net_60967;
  assign seg_16_5_sp4_v_b_36_61079 = net_61079;
  assign seg_16_5_sp4_v_b_42_61085 = net_61085;
  assign seg_16_6_neigh_op_bot_5_60937 = seg_16_5_lutff_5_out_60937;
  assign seg_16_6_sp4_h_r_20_61201 = net_61201;
  assign seg_16_6_sp4_h_r_24_57360 = net_57360;
  assign seg_16_6_sp4_h_r_28_57366 = net_57366;
  assign seg_16_6_sp4_h_r_3_65026 = seg_17_6_sp4_h_r_14_65026;
  assign seg_16_6_sp4_r_v_b_11_64674 = seg_16_4_sp4_r_v_b_35_64674;
  assign seg_16_6_sp4_r_v_b_17_64792 = seg_16_4_sp4_r_v_b_41_64792;
  assign seg_16_6_sp4_r_v_b_21_64796 = seg_16_4_sp4_r_v_b_45_64796;
  assign seg_16_6_sp4_r_v_b_23_64798 = net_64798;
  assign seg_16_6_sp4_r_v_b_35_64920 = net_64920;
  assign seg_16_6_sp4_r_v_b_3_64666 = seg_16_4_sp4_r_v_b_27_64666;
  assign seg_16_6_sp4_v_b_0_60834 = seg_15_5_sp4_r_v_b_13_60834;
  assign seg_16_6_sp4_v_b_10_60844 = seg_15_5_sp4_r_v_b_23_60844;
  assign seg_16_6_sp4_v_b_12_60956 = seg_16_4_sp4_v_b_36_60956;
  assign seg_16_6_sp4_v_b_14_60958 = seg_16_4_sp4_v_b_38_60958;
  assign seg_16_6_sp4_v_b_1_60833 = seg_16_3_sp4_v_b_36_60833;
  assign seg_16_6_sp4_v_b_22_60966 = seg_16_4_sp4_v_b_46_60966;
  assign seg_16_6_sp4_v_b_3_60835 = seg_16_3_sp4_v_b_38_60835;
  assign seg_16_6_sp4_v_b_42_61208 = net_61208;
  assign seg_16_6_sp4_v_b_46_61212 = net_61212;
  assign seg_16_6_sp4_v_b_5_60837 = seg_15_4_sp4_r_v_b_29_60837;
  assign seg_16_6_sp4_v_b_8_60842 = seg_15_5_sp4_r_v_b_21_60842;
  assign seg_16_6_sp4_v_t_36_61325 = seg_16_9_sp4_v_b_12_61325;
  assign seg_16_6_sp4_v_t_46_61335 = seg_15_8_sp4_r_v_b_35_61335;
  assign seg_16_7_lutff_3_out_61181 = net_61181;
  assign seg_16_7_lutff_4_out_61182 = net_61182;
  assign seg_16_7_neigh_op_bnr_4_64890 = seg_17_6_lutff_4_out_64890;
  assign seg_16_7_sp4_h_l_38_49827 = seg_13_7_sp4_h_r_14_49827;
  assign seg_16_7_sp4_h_r_0_65144 = net_65144;
  assign seg_16_7_sp4_h_r_20_61324 = net_61324;
  assign seg_16_7_sp4_h_r_22_61316 = net_61316;
  assign seg_16_7_sp4_h_r_2_65148 = net_65148;
  assign seg_16_7_sp4_h_r_30_57491 = net_57491;
  assign seg_16_7_sp4_h_r_4_65150 = seg_18_7_sp4_h_r_28_65150;
  assign seg_16_7_sp4_r_v_b_13_64911 = net_64911;
  assign seg_16_7_sp4_r_v_b_15_64913 = seg_16_5_sp4_r_v_b_39_64913;
  assign seg_16_7_sp4_r_v_b_29_65037 = net_65037;
  assign seg_16_7_sp4_r_v_b_45_65165 = net_65165;
  assign seg_16_7_sp4_v_b_10_60967 = seg_16_5_sp4_v_b_34_60967;
  assign seg_16_7_sp4_v_b_12_61079 = seg_16_5_sp4_v_b_36_61079;
  assign seg_16_7_sp4_v_b_26_61205 = net_61205;
  assign seg_16_7_sp4_v_b_2_60959 = seg_15_4_sp4_r_v_b_39_60959;
  assign seg_16_7_sp4_v_b_4_60961 = seg_15_4_sp4_r_v_b_41_60961;
  assign seg_16_7_sp4_v_b_5_60960 = seg_15_5_sp4_r_v_b_29_60960;
  assign seg_16_7_sp4_v_b_8_60965 = seg_16_5_sp4_v_b_32_60965;
  assign seg_16_7_sp4_v_b_9_60964 = seg_15_5_sp4_r_v_b_33_60964;
  assign seg_16_8_lutff_0_out_61301 = net_61301;
  assign seg_16_8_sp12_h_r_3_61432 = seg_21_8_sp12_h_r_12_61432;
  assign seg_16_8_sp12_h_r_5_57603 = seg_21_8_sp12_h_r_14_57603;
  assign seg_16_8_sp4_h_l_37_49945 = seg_12_8_sp4_h_r_0_49945;
  assign seg_16_8_sp4_h_l_45_49955 = seg_12_8_sp4_h_r_8_49955;
  assign seg_16_8_sp4_h_r_8_65277 = seg_18_8_sp4_h_r_32_65277;
  assign seg_16_8_sp4_v_b_34_61336 = net_61336;
  assign seg_16_8_sp4_v_b_40_61452 = net_61452;
  assign seg_16_8_sp4_v_b_7_61085 = seg_16_5_sp4_v_b_42_61085;
  assign seg_16_8_sp4_v_t_36_61571 = seg_16_11_sp4_v_b_12_61571;
  assign seg_16_8_sp4_v_t_38_61573 = seg_16_11_sp4_v_b_14_61573;
  assign seg_16_8_sp4_v_t_39_61574 = seg_15_9_sp4_r_v_b_39_61574;
  assign seg_16_8_sp4_v_t_43_61578 = seg_16_12_sp4_v_b_6_61578;
  assign seg_16_9_lutff_4_out_61428 = net_61428;
  assign seg_16_9_lutff_7_out_61431 = net_61431;
  assign seg_16_9_neigh_op_rgt_7_65262 = seg_17_9_lutff_7_out_65262;
  assign seg_16_9_sp12_h_r_12_42402 = net_42402;
  assign seg_16_9_sp4_h_r_24_57729 = net_57729;
  assign seg_16_9_sp4_h_r_34_57731 = net_57731;
  assign seg_16_9_sp4_h_r_42_53908 = net_53908;
  assign seg_16_9_sp4_h_r_46_53902 = net_53902;
  assign seg_16_9_sp4_r_v_b_25_65279 = net_65279;
  assign seg_16_9_sp4_v_b_10_61213 = seg_15_8_sp4_r_v_b_23_61213;
  assign seg_16_9_sp4_v_b_11_61212 = seg_16_6_sp4_v_b_46_61212;
  assign seg_16_9_sp4_v_b_12_61325 = net_61325;
  assign seg_16_9_sp4_v_b_2_61205 = seg_16_7_sp4_v_b_26_61205;
  assign seg_16_9_sp4_v_b_34_61459 = net_61459;
  assign seg_16_9_sp4_v_b_3_61204 = seg_15_9_sp4_r_v_b_3_61204;
  assign seg_16_9_sp4_v_b_42_61577 = net_61577;
  assign seg_16_9_sp4_v_b_7_61208 = seg_16_6_sp4_v_b_42_61208;
  assign seg_17_0_span4_horz_r_12_56601 = net_56601;
  assign seg_17_0_span4_vert_32_64408 = net_64408;
  assign seg_17_10_lutff_0_out_65378 = net_65378;
  assign seg_17_10_lutff_1_out_65379 = net_65379;
  assign seg_17_10_lutff_2_out_65380 = net_65380;
  assign seg_17_10_lutff_5_out_65383 = net_65383;
  assign seg_17_10_lutff_7_out_65385 = net_65385;
  assign seg_17_10_neigh_op_rgt_3_69212 = seg_18_10_lutff_3_out_69212;
  assign seg_17_10_neigh_op_rgt_6_69215 = seg_18_10_lutff_6_out_69215;
  assign seg_17_10_sp12_h_r_14_42526 = net_42526;
  assign seg_17_10_sp4_h_l_38_54027 = seg_14_10_sp4_h_r_14_54027;
  assign seg_17_10_sp4_h_l_40_54029 = seg_14_10_sp4_h_r_16_54029;
  assign seg_17_10_sp4_h_l_42_54031 = seg_14_10_sp4_h_r_18_54031;
  assign seg_17_10_sp4_h_l_43_54030 = seg_15_10_sp4_h_r_30_54030;
  assign seg_17_10_sp4_h_l_44_54033 = seg_14_10_sp4_h_r_20_54033;
  assign seg_17_10_sp4_h_l_46_54025 = seg_14_10_sp4_h_r_22_54025;
  assign seg_17_10_sp4_h_r_24_61682 = net_61682;
  assign seg_17_10_sp4_h_r_26_61686 = net_61686;
  assign seg_17_10_sp4_r_v_b_11_68997 = net_68997;
  assign seg_17_10_sp4_v_b_10_65167 = net_65167;
  assign seg_17_10_sp4_v_b_26_65405 = net_65405;
  assign seg_17_10_sp4_v_b_8_65165 = seg_16_7_sp4_r_v_b_45_65165;
  assign seg_17_11_lutff_1_out_65502 = net_65502;
  assign seg_17_11_lutff_2_out_65503 = net_65503;
  assign seg_17_11_lutff_3_out_65504 = net_65504;
  assign seg_17_11_lutff_4_out_65505 = net_65505;
  assign seg_17_11_lutff_5_out_65506 = net_65506;
  assign seg_17_11_lutff_6_out_65507 = net_65507;
  assign seg_17_11_lutff_7_out_65508 = net_65508;
  assign seg_17_11_neigh_op_bot_0_65378 = seg_17_10_lutff_0_out_65378;
  assign seg_17_11_neigh_op_bot_1_65379 = seg_17_10_lutff_1_out_65379;
  assign seg_17_11_neigh_op_bot_5_65383 = seg_17_10_lutff_5_out_65383;
  assign seg_17_11_neigh_op_lft_5_61675 = seg_16_11_lutff_5_out_61675;
  assign seg_17_11_neigh_op_rgt_0_69332 = seg_18_11_lutff_0_out_69332;
  assign seg_17_11_neigh_op_rgt_2_69334 = seg_18_11_lutff_2_out_69334;
  assign seg_17_11_neigh_op_tnr_0_69455 = seg_18_12_lutff_0_out_69455;
  assign seg_17_11_neigh_op_tnr_2_69457 = seg_18_12_lutff_2_out_69457;
  assign seg_17_11_neigh_op_tnr_6_69461 = seg_18_12_lutff_6_out_69461;
  assign seg_17_11_neigh_op_top_0_65624 = seg_17_12_lutff_0_out_65624;
  assign seg_17_11_neigh_op_top_4_65628 = seg_17_12_lutff_4_out_65628;
  assign seg_17_11_neigh_op_top_7_65631 = seg_17_12_lutff_7_out_65631;
  assign seg_17_11_sp12_v_b_14_68850 = net_68850;
  assign seg_17_11_sp4_h_l_36_54146 = seg_16_11_sp4_h_r_36_54146;
  assign seg_17_11_sp4_h_l_45_54155 = seg_13_11_sp4_h_r_8_54155;
  assign seg_17_11_sp4_h_r_46_57978 = seg_15_11_sp4_h_r_22_57978;
  assign seg_17_11_sp4_v_b_10_65290 = seg_16_10_sp4_r_v_b_23_65290;
  assign seg_17_11_sp4_v_b_12_65402 = net_65402;
  assign seg_17_11_sp4_v_b_1_65279 = seg_16_9_sp4_r_v_b_25_65279;
  assign seg_17_11_sp4_v_b_4_65284 = seg_16_10_sp4_r_v_b_17_65284;
  assign seg_17_11_sp4_v_b_8_65288 = seg_16_10_sp4_r_v_b_21_65288;
  assign seg_17_11_sp4_v_t_42_65777 = seg_16_13_sp4_r_v_b_31_65777;
  assign seg_17_12_lutff_0_out_65624 = net_65624;
  assign seg_17_12_lutff_1_out_65625 = net_65625;
  assign seg_17_12_lutff_2_out_65626 = net_65626;
  assign seg_17_12_lutff_3_out_65627 = net_65627;
  assign seg_17_12_lutff_4_out_65628 = net_65628;
  assign seg_17_12_lutff_5_out_65629 = net_65629;
  assign seg_17_12_lutff_6_out_65630 = net_65630;
  assign seg_17_12_lutff_7_out_65631 = net_65631;
  assign seg_17_12_neigh_op_bnl_1_61671 = seg_16_11_lutff_1_out_61671;
  assign seg_17_12_neigh_op_bnl_3_61673 = seg_16_11_lutff_3_out_61673;
  assign seg_17_12_sp4_v_b_46_65781 = seg_16_15_sp4_r_v_b_11_65781;
  assign seg_17_12_sp4_v_b_5_65406 = seg_16_10_sp4_r_v_b_29_65406;
  assign seg_17_12_sp4_v_b_7_65408 = seg_16_10_sp4_r_v_b_31_65408;
  assign seg_17_12_sp4_v_b_8_65411 = seg_16_11_sp4_r_v_b_21_65411;
  assign seg_17_12_sp4_v_b_9_65410 = seg_16_10_sp4_r_v_b_33_65410;
  assign seg_17_12_sp4_v_t_36_65894 = seg_17_15_sp4_v_b_12_65894;
  assign seg_17_13_lutff_2_out_65749 = net_65749;
  assign seg_17_13_lutff_3_out_65750 = net_65750;
  assign seg_17_13_lutff_4_out_65751 = net_65751;
  assign seg_17_13_lutff_5_out_65752 = net_65752;
  assign seg_17_13_lutff_6_out_65753 = net_65753;
  assign seg_17_13_neigh_op_tnl_1_62040 = seg_16_14_lutff_1_out_62040;
  assign seg_17_13_neigh_op_tnl_2_62041 = seg_16_14_lutff_2_out_62041;
  assign seg_17_13_neigh_op_tnl_3_62042 = seg_16_14_lutff_3_out_62042;
  assign seg_17_13_neigh_op_tnl_4_62043 = seg_16_14_lutff_4_out_62043;
  assign seg_17_13_neigh_op_tnl_5_62044 = seg_16_14_lutff_5_out_62044;
  assign seg_17_13_neigh_op_tnl_6_62045 = seg_16_14_lutff_6_out_62045;
  assign seg_17_13_neigh_op_tnl_7_62046 = seg_16_14_lutff_7_out_62046;
  assign seg_17_13_neigh_op_top_4_65874 = seg_17_14_lutff_4_out_65874;
  assign seg_17_13_sp4_h_r_2_69717 = net_69717;
  assign seg_17_13_sp4_v_b_2_65528 = seg_16_10_sp4_r_v_b_39_65528;
  assign seg_17_13_sp4_v_b_4_65530 = seg_16_10_sp4_r_v_b_41_65530;
  assign seg_17_13_sp4_v_b_6_65532 = seg_16_10_sp4_r_v_b_43_65532;
  assign seg_17_14_lutff_1_out_65871 = net_65871;
  assign seg_17_14_lutff_2_out_65872 = net_65872;
  assign seg_17_14_lutff_3_out_65873 = net_65873;
  assign seg_17_14_lutff_4_out_65874 = net_65874;
  assign seg_17_14_lutff_5_out_65875 = net_65875;
  assign seg_17_14_lutff_6_out_65876 = net_65876;
  assign seg_17_14_lutff_7_out_65877 = net_65877;
  assign seg_17_14_neigh_op_bot_2_65749 = seg_17_13_lutff_2_out_65749;
  assign seg_17_14_neigh_op_bot_3_65750 = seg_17_13_lutff_3_out_65750;
  assign seg_17_14_neigh_op_bot_4_65751 = seg_17_13_lutff_4_out_65751;
  assign seg_17_14_neigh_op_bot_5_65752 = seg_17_13_lutff_5_out_65752;
  assign seg_17_14_neigh_op_bot_6_65753 = seg_17_13_lutff_6_out_65753;
  assign seg_17_14_neigh_op_tnl_0_62162 = seg_16_15_lutff_0_out_62162;
  assign seg_17_14_neigh_op_top_4_65997 = seg_17_15_lutff_4_out_65997;
  assign seg_17_14_neigh_op_top_7_66000 = seg_17_15_lutff_7_out_66000;
  assign seg_17_14_sp4_h_l_39_54518 = seg_13_14_sp4_h_r_2_54518;
  assign seg_17_14_sp4_h_r_0_69836 = net_69836;
  assign seg_17_14_sp4_h_r_3_69841 = seg_20_14_sp4_h_r_38_69841;
  assign seg_17_14_sp4_v_b_28_65899 = seg_17_16_sp4_v_b_4_65899;
  assign seg_17_14_sp4_v_b_2_65651 = seg_16_13_sp4_r_v_b_15_65651;
  assign seg_17_14_sp4_v_b_30_65901 = seg_17_16_sp4_v_b_6_65901;
  assign seg_17_14_sp4_v_b_32_65903 = seg_17_16_sp4_v_b_8_65903;
  assign seg_17_14_sp4_v_b_34_65905 = seg_17_16_sp4_v_b_10_65905;
  assign seg_17_14_sp4_v_b_36_66017 = seg_17_16_sp4_v_b_12_66017;
  assign seg_17_14_sp4_v_b_40_66021 = net_66021;
  assign seg_17_14_sp4_v_t_38_66142 = seg_17_17_sp4_v_b_14_66142;
  assign seg_17_15_lutff_0_out_65993 = net_65993;
  assign seg_17_15_lutff_1_out_65994 = net_65994;
  assign seg_17_15_lutff_2_out_65995 = net_65995;
  assign seg_17_15_lutff_3_out_65996 = net_65996;
  assign seg_17_15_lutff_4_out_65997 = net_65997;
  assign seg_17_15_lutff_5_out_65998 = net_65998;
  assign seg_17_15_lutff_6_out_65999 = net_65999;
  assign seg_17_15_lutff_7_out_66000 = net_66000;
  assign seg_17_15_neigh_op_tnl_2_62287 = seg_16_16_lutff_2_out_62287;
  assign seg_17_15_neigh_op_tnl_3_62288 = seg_16_16_lutff_3_out_62288;
  assign seg_17_15_neigh_op_tnr_2_69949 = seg_18_16_lutff_2_out_69949;
  assign seg_17_15_neigh_op_tnr_5_69952 = seg_18_16_lutff_5_out_69952;
  assign seg_17_15_sp4_h_r_4_69965 = net_69965;
  assign seg_17_15_sp4_r_v_b_27_69850 = seg_17_17_sp4_r_v_b_3_69850;
  assign seg_17_15_sp4_r_v_b_3_69604 = net_69604;
  assign seg_17_15_sp4_r_v_b_9_69610 = net_69610;
  assign seg_17_15_sp4_v_b_12_65894 = net_65894;
  assign seg_17_15_sp4_v_b_27_66019 = seg_16_17_sp4_r_v_b_3_66019;
  assign seg_17_15_sp4_v_b_33_66025 = seg_16_17_sp4_r_v_b_9_66025;
  assign seg_17_15_sp4_v_b_37_66141 = seg_16_17_sp4_r_v_b_13_66141;
  assign seg_17_15_sp4_v_b_7_65777 = seg_16_13_sp4_r_v_b_31_65777;
  assign seg_17_16_lutff_1_out_66117 = net_66117;
  assign seg_17_16_neigh_op_bnr_1_69825 = seg_18_15_lutff_1_out_69825;
  assign seg_17_16_neigh_op_bnr_2_69826 = seg_18_15_lutff_2_out_69826;
  assign seg_17_16_neigh_op_bnr_3_69827 = seg_18_15_lutff_3_out_69827;
  assign seg_17_16_neigh_op_bnr_4_69828 = seg_18_15_lutff_4_out_69828;
  assign seg_17_16_neigh_op_bnr_5_69829 = seg_18_15_lutff_5_out_69829;
  assign seg_17_16_neigh_op_bnr_6_69830 = seg_18_15_lutff_6_out_69830;
  assign seg_17_16_neigh_op_bnr_7_69831 = seg_18_15_lutff_7_out_69831;
  assign seg_17_16_neigh_op_rgt_4_69951 = seg_18_16_lutff_4_out_69951;
  assign seg_17_16_neigh_op_tnr_4_70074 = seg_18_17_lutff_4_out_70074;
  assign seg_17_16_sp4_v_b_10_65905 = net_65905;
  assign seg_17_16_sp4_v_b_11_65904 = seg_16_16_sp4_r_v_b_11_65904;
  assign seg_17_16_sp4_v_b_12_66017 = net_66017;
  assign seg_17_16_sp4_v_b_4_65899 = net_65899;
  assign seg_17_16_sp4_v_b_6_65901 = net_65901;
  assign seg_17_16_sp4_v_b_8_65903 = net_65903;
  assign seg_17_16_sp4_v_t_41_66391 = seg_17_18_sp4_v_b_28_66391;
  assign seg_17_16_sp4_v_t_43_66393 = seg_16_17_sp4_r_v_b_43_66393;
  assign seg_17_17_lutff_0_out_66239 = net_66239;
  assign seg_17_17_lutff_3_out_66242 = net_66242;
  assign seg_17_17_lutff_4_out_66243 = net_66243;
  assign seg_17_17_lutff_5_out_66244 = net_66244;
  assign seg_17_17_neigh_op_bnr_0_69947 = seg_18_16_lutff_0_out_69947;
  assign seg_17_17_neigh_op_bnr_4_69951 = seg_18_16_lutff_4_out_69951;
  assign seg_17_17_neigh_op_bot_1_66117 = seg_17_16_lutff_1_out_66117;
  assign seg_17_17_neigh_op_rgt_4_70074 = seg_18_17_lutff_4_out_70074;
  assign seg_17_17_neigh_op_top_6_66368 = seg_17_18_lutff_6_out_66368;
  assign seg_17_17_sp4_h_r_14_66379 = net_66379;
  assign seg_17_17_sp4_h_r_24_62543 = net_62543;
  assign seg_17_17_sp4_h_r_39_58717 = seg_14_17_sp4_h_r_2_58717;
  assign seg_17_17_sp4_h_r_40_58720 = net_58720;
  assign seg_17_17_sp4_h_r_46_58716 = net_58716;
  assign seg_17_17_sp4_r_v_b_13_69972 = net_69972;
  assign seg_17_17_sp4_r_v_b_3_69850 = net_69850;
  assign seg_17_17_sp4_v_b_14_66142 = net_66142;
  assign seg_17_17_sp4_v_b_5_66021 = seg_17_14_sp4_v_b_40_66021;
  assign seg_17_18_lutff_6_out_66368 = net_66368;
  assign seg_17_18_neigh_op_bot_4_66243 = seg_17_17_lutff_4_out_66243;
  assign seg_17_18_sp12_v_b_1_68850 = seg_17_11_sp12_v_b_14_68850;
  assign seg_17_18_sp4_h_r_44_58847 = net_58847;
  assign seg_17_18_sp4_v_b_28_66391 = net_66391;
  assign seg_17_2_sp4_h_r_0_68360 = net_68360;
  assign seg_17_2_sp4_h_r_14_64534 = net_64534;
  assign seg_17_3_lutff_0_out_64517 = net_64517;
  assign seg_17_3_lutff_1_out_64518 = net_64518;
  assign seg_17_3_lutff_3_out_64520 = net_64520;
  assign seg_17_3_lutff_4_out_64521 = net_64521;
  assign seg_17_3_sp4_h_l_39_53165 = seg_13_3_sp4_h_r_2_53165;
  assign seg_17_3_sp4_h_l_47_53163 = seg_13_3_sp4_h_r_10_53163;
  assign seg_17_3_sp4_h_r_11_68486 = seg_20_3_sp4_h_r_46_68486;
  assign seg_17_3_sp4_h_r_36_56992 = net_56992;
  assign seg_17_3_sp4_h_r_3_68488 = seg_20_3_sp4_h_r_38_68488;
  assign seg_17_3_sp4_v_b_8_64408 = seg_17_0_span4_vert_32_64408;
  assign seg_17_4_lutff_0_out_64640 = net_64640;
  assign seg_17_4_lutff_1_out_64641 = net_64641;
  assign seg_17_4_lutff_3_out_64643 = net_64643;
  assign seg_17_4_lutff_4_out_64644 = net_64644;
  assign seg_17_4_lutff_5_out_64645 = net_64645;
  assign seg_17_4_lutff_6_out_64646 = net_64646;
  assign seg_17_4_lutff_7_out_64647 = net_64647;
  assign seg_17_4_sp12_h_r_3_64771 = seg_22_4_sp12_h_r_12_64771;
  assign seg_17_4_sp4_h_l_37_53284 = seg_15_4_sp4_h_r_24_53284;
  assign seg_17_4_sp4_h_l_39_53288 = seg_15_4_sp4_h_r_26_53288;
  assign seg_17_4_sp4_h_l_44_53295 = seg_14_4_sp4_h_r_20_53295;
  assign seg_17_4_sp4_h_l_47_53286 = seg_15_4_sp4_h_r_34_53286;
  assign seg_17_4_sp4_r_v_b_32_68504 = seg_18_6_sp4_v_b_8_68504;
  assign seg_17_4_sp4_r_v_b_5_68248 = net_68248;
  assign seg_17_4_sp4_v_b_10_64424 = seg_16_3_sp4_r_v_b_23_64424;
  assign seg_17_4_sp4_v_t_38_64912 = seg_17_7_sp4_v_b_14_64912;
  assign seg_17_5_lutff_0_out_64763 = net_64763;
  assign seg_17_5_lutff_1_out_64764 = net_64764;
  assign seg_17_5_lutff_2_out_64765 = net_64765;
  assign seg_17_5_lutff_3_out_64766 = net_64766;
  assign seg_17_5_lutff_5_out_64768 = net_64768;
  assign seg_17_5_lutff_6_out_64769 = net_64769;
  assign seg_17_5_lutff_7_out_64770 = net_64770;
  assign seg_17_5_sp4_h_l_37_53407 = seg_15_5_sp4_h_r_24_53407;
  assign seg_17_5_sp4_h_l_39_53411 = seg_15_5_sp4_h_r_26_53411;
  assign seg_17_5_sp4_h_l_43_53415 = seg_15_5_sp4_h_r_30_53415;
  assign seg_17_5_sp4_h_r_11_68732 = seg_20_5_sp4_h_r_46_68732;
  assign seg_17_5_sp4_h_r_1_68730 = seg_20_5_sp4_h_r_36_68730;
  assign seg_17_5_sp4_h_r_3_68734 = seg_20_5_sp4_h_r_38_68734;
  assign seg_17_5_sp4_h_r_5_68736 = seg_20_5_sp4_h_r_40_68736;
  assign seg_17_5_sp4_h_r_7_68738 = seg_20_5_sp4_h_r_42_68738;
  assign seg_17_5_sp4_r_v_b_47_68752 = seg_18_8_sp4_v_b_10_68752;
  assign seg_17_5_sp4_v_t_45_65042 = seg_17_9_sp4_v_b_8_65042;
  assign seg_17_6_lutff_2_out_64888 = net_64888;
  assign seg_17_6_lutff_4_out_64890 = net_64890;
  assign seg_17_6_lutff_5_out_64891 = net_64891;
  assign seg_17_6_lutff_6_out_64892 = net_64892;
  assign seg_17_6_neigh_op_rgt_3_68720 = seg_18_6_lutff_3_out_68720;
  assign seg_17_6_sp4_h_l_37_53530 = seg_13_6_sp4_h_r_0_53530;
  assign seg_17_6_sp4_h_l_47_53532 = seg_13_6_sp4_h_r_10_53532;
  assign seg_17_6_sp4_h_r_14_65026 = net_65026;
  assign seg_17_6_sp4_h_r_5_68859 = seg_20_6_sp4_h_r_40_68859;
  assign seg_17_6_sp4_v_b_0_64665 = seg_16_3_sp4_r_v_b_37_64665;
  assign seg_17_6_sp4_v_t_47_65167 = seg_17_10_sp4_v_b_10_65167;
  assign seg_17_7_lutff_7_out_65016 = net_65016;
  assign seg_17_7_sp4_h_r_3_68980 = seg_18_7_sp4_h_r_14_68980;
  assign seg_17_7_sp4_h_r_46_57486 = net_57486;
  assign seg_17_7_sp4_h_r_7_68984 = seg_20_7_sp4_h_r_42_68984;
  assign seg_17_7_sp4_h_r_9_68986 = seg_18_7_sp4_h_r_20_68986;
  assign seg_17_7_sp4_v_b_10_64798 = seg_16_6_sp4_r_v_b_23_64798;
  assign seg_17_7_sp4_v_b_14_64912 = net_64912;
  assign seg_17_8_sp4_h_l_36_53777 = seg_14_8_sp4_h_r_12_53777;
  assign seg_17_8_sp4_h_l_39_53780 = seg_13_8_sp4_h_r_2_53780;
  assign seg_17_8_sp4_h_l_47_53778 = seg_15_8_sp4_h_r_34_53778;
  assign seg_17_8_sp4_h_r_34_61438 = net_61438;
  assign seg_17_8_sp4_h_r_36_57607 = net_57607;
  assign seg_17_8_sp4_h_r_44_57617 = net_57617;
  assign seg_17_8_sp4_h_r_7_69107 = seg_18_8_sp4_h_r_18_69107;
  assign seg_17_8_sp4_v_b_0_64911 = seg_16_7_sp4_r_v_b_13_64911;
  assign seg_17_8_sp4_v_b_11_64920 = seg_16_6_sp4_r_v_b_35_64920;
  assign seg_17_8_sp4_v_t_36_65402 = seg_17_11_sp4_v_b_12_65402;
  assign seg_17_8_sp4_v_t_39_65405 = seg_17_10_sp4_v_b_26_65405;
  assign seg_17_9_lutff_7_out_65262 = net_65262;
  assign seg_17_9_sp4_h_l_41_53905 = seg_15_9_sp4_h_r_28_53905;
  assign seg_17_9_sp4_h_l_45_53909 = seg_15_9_sp4_h_r_32_53909;
  assign seg_17_9_sp4_h_r_7_69230 = seg_20_9_sp4_h_r_42_69230;
  assign seg_17_9_sp4_v_b_5_65037 = seg_16_7_sp4_r_v_b_29_65037;
  assign seg_17_9_sp4_v_b_8_65042 = net_65042;
  assign seg_18_0_span4_horz_r_12_60431 = net_60431;
  assign seg_18_10_lutff_1_out_69210 = net_69210;
  assign seg_18_10_lutff_3_out_69212 = net_69212;
  assign seg_18_10_lutff_4_out_69213 = net_69213;
  assign seg_18_10_lutff_6_out_69215 = net_69215;
  assign seg_18_10_neigh_op_bot_5_69091 = seg_18_9_lutff_5_out_69091;
  assign seg_18_10_neigh_op_bot_6_69092 = seg_18_9_lutff_6_out_69092;
  assign seg_18_10_neigh_op_lft_2_65380 = seg_17_10_lutff_2_out_65380;
  assign seg_18_10_neigh_op_top_7_69339 = seg_18_11_lutff_7_out_69339;
  assign seg_18_10_sp4_h_r_0_73175 = seg_20_10_sp4_h_r_24_73175;
  assign seg_18_10_sp4_h_r_26_65517 = net_65517;
  assign seg_18_10_sp4_h_r_30_65521 = net_65521;
  assign seg_18_10_sp4_h_r_5_73182 = seg_21_10_sp4_h_r_40_73182;
  assign seg_18_10_sp4_r_v_b_21_72950 = net_72950;
  assign seg_18_10_sp4_v_b_1_68987 = seg_18_7_sp4_v_b_36_68987;
  assign seg_18_10_sp4_v_b_38_69358 = seg_18_12_sp4_v_b_14_69358;
  assign seg_18_10_sp4_v_b_3_68989 = seg_18_7_sp4_v_b_38_68989;
  assign seg_18_10_sp4_v_b_47_69367 = seg_18_13_sp4_v_b_10_69367;
  assign seg_18_10_sp4_v_b_7_68993 = seg_18_7_sp4_v_b_42_68993;
  assign seg_18_10_sp4_v_b_8_68996 = seg_18_8_sp4_v_b_32_68996;
  assign seg_18_10_sp4_v_b_9_68995 = seg_18_7_sp4_v_b_44_68995;
  assign seg_18_11_lutff_0_out_69332 = net_69332;
  assign seg_18_11_lutff_1_out_69333 = net_69333;
  assign seg_18_11_lutff_2_out_69334 = net_69334;
  assign seg_18_11_lutff_3_out_69335 = net_69335;
  assign seg_18_11_lutff_5_out_69337 = net_69337;
  assign seg_18_11_lutff_6_out_69338 = net_69338;
  assign seg_18_11_lutff_7_out_69339 = net_69339;
  assign seg_18_11_neigh_op_lft_6_65507 = seg_17_11_lutff_6_out_65507;
  assign seg_18_11_neigh_op_lft_7_65508 = seg_17_11_lutff_7_out_65508;
  assign seg_18_11_sp4_h_l_37_57975 = seg_16_11_sp4_h_r_24_57975;
  assign seg_18_11_sp4_h_r_24_65636 = net_65636;
  assign seg_18_11_sp4_h_r_32_65646 = seg_16_11_sp4_h_r_8_65646;
  assign seg_18_11_sp4_h_r_40_61812 = net_61812;
  assign seg_18_11_sp4_h_r_6_73306 = seg_20_11_sp4_h_r_30_73306;
  assign seg_18_11_sp4_h_r_8_73308 = net_73308;
  assign seg_18_11_sp4_v_b_24_69357 = net_69357;
  assign seg_18_11_sp4_v_t_36_69602 = seg_18_14_sp4_v_b_12_69602;
  assign seg_18_12_lutff_0_out_69455 = net_69455;
  assign seg_18_12_lutff_1_out_69456 = net_69456;
  assign seg_18_12_lutff_2_out_69457 = net_69457;
  assign seg_18_12_lutff_3_out_69458 = net_69458;
  assign seg_18_12_lutff_4_out_69459 = net_69459;
  assign seg_18_12_lutff_6_out_69461 = net_69461;
  assign seg_18_12_neigh_op_lft_1_65625 = seg_17_12_lutff_1_out_65625;
  assign seg_18_12_neigh_op_top_0_69578 = seg_18_13_lutff_0_out_69578;
  assign seg_18_12_sp4_v_b_14_69358 = net_69358;
  assign seg_18_12_sp4_v_t_39_69728 = seg_18_16_sp4_v_b_2_69728;
  assign seg_18_13_lutff_0_out_69578 = net_69578;
  assign seg_18_13_neigh_op_top_1_69702 = seg_18_14_lutff_1_out_69702;
  assign seg_18_13_sp4_h_r_34_65884 = net_65884;
  assign seg_18_13_sp4_h_r_36_62052 = net_62052;
  assign seg_18_13_sp4_h_r_40_62058 = net_62058;
  assign seg_18_13_sp4_h_r_44_62062 = net_62062;
  assign seg_18_13_sp4_v_b_0_69357 = seg_18_11_sp4_v_b_24_69357;
  assign seg_18_13_sp4_v_b_10_69367 = net_69367;
  assign seg_18_13_sp4_v_b_27_69604 = seg_17_15_sp4_r_v_b_3_69604;
  assign seg_18_13_sp4_v_b_33_69610 = seg_17_15_sp4_r_v_b_9_69610;
  assign seg_18_13_sp4_v_b_41_69730 = seg_18_16_sp4_v_b_4_69730;
  assign seg_18_13_sp4_v_b_47_69736 = seg_18_16_sp4_v_b_10_69736;
  assign seg_18_14_lutff_0_out_69701 = net_69701;
  assign seg_18_14_lutff_1_out_69702 = net_69702;
  assign seg_18_14_lutff_2_out_69703 = net_69703;
  assign seg_18_14_lutff_3_out_69704 = net_69704;
  assign seg_18_14_lutff_4_out_69705 = net_69705;
  assign seg_18_14_lutff_7_out_69708 = net_69708;
  assign seg_18_14_neigh_op_lft_1_65871 = seg_17_14_lutff_1_out_65871;
  assign seg_18_14_neigh_op_lft_2_65872 = seg_17_14_lutff_2_out_65872;
  assign seg_18_14_neigh_op_lft_3_65873 = seg_17_14_lutff_3_out_65873;
  assign seg_18_14_neigh_op_lft_6_65876 = seg_17_14_lutff_6_out_65876;
  assign seg_18_14_sp4_h_l_41_58350 = seg_14_14_sp4_h_r_4_58350;
  assign seg_18_14_sp4_h_l_44_58355 = seg_15_14_sp4_h_r_20_58355;
  assign seg_18_14_sp4_h_l_45_58354 = seg_14_14_sp4_h_r_8_58354;
  assign seg_18_14_sp4_h_l_47_58346 = seg_14_14_sp4_h_r_10_58346;
  assign seg_18_14_sp4_h_r_30_66013 = net_66013;
  assign seg_18_14_sp4_h_r_32_66015 = net_66015;
  assign seg_18_14_sp4_h_r_36_62175 = net_62175;
  assign seg_18_14_sp4_h_r_38_62179 = net_62179;
  assign seg_18_14_sp4_h_r_40_62181 = net_62181;
  assign seg_18_14_sp4_h_r_41_62180 = seg_15_14_sp4_h_r_4_62180;
  assign seg_18_14_sp4_r_v_b_11_73320 = net_73320;
  assign seg_18_14_sp4_v_b_12_69602 = net_69602;
  assign seg_18_14_sp4_v_t_37_69972 = seg_17_17_sp4_r_v_b_13_69972;
  assign seg_18_14_sp4_v_t_43_69978 = seg_18_16_sp4_v_b_30_69978;
  assign seg_18_15_lutff_1_out_69825 = net_69825;
  assign seg_18_15_lutff_2_out_69826 = net_69826;
  assign seg_18_15_lutff_3_out_69827 = net_69827;
  assign seg_18_15_lutff_4_out_69828 = net_69828;
  assign seg_18_15_lutff_5_out_69829 = net_69829;
  assign seg_18_15_lutff_6_out_69830 = net_69830;
  assign seg_18_15_lutff_7_out_69831 = net_69831;
  assign seg_18_15_neigh_op_bot_0_69701 = seg_18_14_lutff_0_out_69701;
  assign seg_18_15_neigh_op_bot_2_69703 = seg_18_14_lutff_2_out_69703;
  assign seg_18_15_neigh_op_bot_3_69704 = seg_18_14_lutff_3_out_69704;
  assign seg_18_15_neigh_op_bot_4_69705 = seg_18_14_lutff_4_out_69705;
  assign seg_18_15_neigh_op_bot_7_69708 = seg_18_14_lutff_7_out_69708;
  assign seg_18_15_neigh_op_lft_1_65994 = seg_17_15_lutff_1_out_65994;
  assign seg_18_15_neigh_op_lft_4_65997 = seg_17_15_lutff_4_out_65997;
  assign seg_18_15_neigh_op_lft_5_65998 = seg_17_15_lutff_5_out_65998;
  assign seg_18_15_neigh_op_lft_6_65999 = seg_17_15_lutff_6_out_65999;
  assign seg_18_15_neigh_op_lft_7_66000 = seg_17_15_lutff_7_out_66000;
  assign seg_18_15_neigh_op_top_2_69949 = seg_18_16_lutff_2_out_69949;
  assign seg_18_15_neigh_op_top_5_69952 = seg_18_16_lutff_5_out_69952;
  assign seg_18_15_sp4_h_l_37_58467 = seg_16_15_sp4_h_r_24_58467;
  assign seg_18_15_sp4_h_r_17_69965 = seg_17_15_sp4_h_r_4_69965;
  assign seg_18_15_sp4_h_r_34_66130 = seg_16_15_sp4_h_r_10_66130;
  assign seg_18_15_sp4_h_r_36_62298 = seg_16_15_sp4_h_r_12_62298;
  assign seg_18_15_sp4_v_b_43_69978 = seg_18_16_sp4_v_b_30_69978;
  assign seg_18_16_lutff_0_out_69947 = net_69947;
  assign seg_18_16_lutff_1_out_69948 = net_69948;
  assign seg_18_16_lutff_2_out_69949 = net_69949;
  assign seg_18_16_lutff_4_out_69951 = net_69951;
  assign seg_18_16_lutff_5_out_69952 = net_69952;
  assign seg_18_16_neigh_op_bnl_4_65997 = seg_17_15_lutff_4_out_65997;
  assign seg_18_16_neigh_op_bnl_7_66000 = seg_17_15_lutff_7_out_66000;
  assign seg_18_16_neigh_op_tnl_0_66239 = seg_17_17_lutff_0_out_66239;
  assign seg_18_16_sp12_v_b_1_72435 = seg_18_7_sp12_v_b_18_72435;
  assign seg_18_16_sp4_h_r_32_66261 = seg_16_16_sp4_h_r_8_66261;
  assign seg_18_16_sp4_h_r_34_66253 = net_66253;
  assign seg_18_16_sp4_v_b_10_69736 = net_69736;
  assign seg_18_16_sp4_v_b_2_69728 = net_69728;
  assign seg_18_16_sp4_v_b_30_69978 = net_69978;
  assign seg_18_16_sp4_v_b_4_69730 = net_69730;
  assign seg_18_17_lutff_4_out_70074 = net_70074;
  assign seg_18_17_sp4_h_r_39_62547 = seg_15_17_sp4_h_r_2_62547;
  assign seg_18_2_sp4_h_r_12_68361 = seg_20_2_sp4_h_r_36_68361;
  assign seg_18_2_sp4_h_r_22_68363 = seg_20_2_sp4_h_r_46_68363;
  assign seg_18_2_sp4_h_r_24_64529 = net_64529;
  assign seg_18_2_sp4_h_r_40_60705 = net_60705;
  assign seg_18_3_lutff_0_out_68348 = net_68348;
  assign seg_18_3_lutff_1_out_68349 = net_68349;
  assign seg_18_3_lutff_2_out_68350 = net_68350;
  assign seg_18_3_lutff_3_out_68351 = net_68351;
  assign seg_18_3_lutff_4_out_68352 = net_68352;
  assign seg_18_3_lutff_5_out_68353 = net_68353;
  assign seg_18_3_lutff_7_out_68355 = net_68355;
  assign seg_18_3_sp4_h_r_11_72317 = seg_21_3_sp4_h_r_46_72317;
  assign seg_18_3_sp4_h_r_18_68492 = seg_20_3_sp4_h_r_42_68492;
  assign seg_18_3_sp4_h_r_1_72315 = seg_21_3_sp4_h_r_36_72315;
  assign seg_18_3_sp4_h_r_4_72320 = seg_20_3_sp4_h_r_28_72320;
  assign seg_18_3_sp4_v_b_44_68503 = net_68503;
  assign seg_18_4_neigh_op_bnl_1_64518 = seg_17_3_lutff_1_out_64518;
  assign seg_18_4_neigh_op_bot_0_68348 = seg_18_3_lutff_0_out_68348;
  assign seg_18_4_neigh_op_bot_1_68349 = seg_18_3_lutff_1_out_68349;
  assign seg_18_4_neigh_op_bot_2_68350 = seg_18_3_lutff_2_out_68350;
  assign seg_18_4_neigh_op_bot_3_68351 = seg_18_3_lutff_3_out_68351;
  assign seg_18_4_neigh_op_bot_4_68352 = seg_18_3_lutff_4_out_68352;
  assign seg_18_4_neigh_op_bot_7_68355 = seg_18_3_lutff_7_out_68355;
  assign seg_18_4_neigh_op_tnl_5_64768 = seg_17_5_lutff_5_out_64768;
  assign seg_18_4_neigh_op_top_2_68596 = seg_18_5_lutff_2_out_68596;
  assign seg_18_4_neigh_op_top_4_68598 = seg_18_5_lutff_4_out_68598;
  assign seg_18_4_neigh_op_top_6_68600 = seg_18_5_lutff_6_out_68600;
  assign seg_18_4_neigh_op_top_7_68601 = seg_18_5_lutff_7_out_68601;
  assign seg_18_4_sp4_h_r_11_72440 = seg_21_4_sp4_h_r_46_72440;
  assign seg_18_4_sp4_h_r_1_72438 = seg_21_4_sp4_h_r_36_72438;
  assign seg_18_4_sp4_h_r_2_72441 = net_72441;
  assign seg_18_4_sp4_h_r_7_72446 = seg_21_4_sp4_h_r_42_72446;
  assign seg_18_4_sp4_r_v_b_45_72458 = net_72458;
  assign seg_18_4_sp4_r_v_b_47_72460 = net_72460;
  assign seg_18_4_sp4_v_b_24_68496 = seg_18_6_sp4_v_b_0_68496;
  assign seg_18_4_sp4_v_b_36_68618 = net_68618;
  assign seg_18_4_sp4_v_b_38_68620 = net_68620;
  assign seg_18_4_sp4_v_b_40_68622 = net_68622;
  assign seg_18_4_sp4_v_b_42_68624 = net_68624;
  assign seg_18_4_sp4_v_b_5_68248 = seg_17_4_sp4_r_v_b_5_68248;
  assign seg_18_5_lutff_2_out_68596 = net_68596;
  assign seg_18_5_lutff_3_out_68597 = net_68597;
  assign seg_18_5_lutff_4_out_68598 = net_68598;
  assign seg_18_5_lutff_5_out_68599 = net_68599;
  assign seg_18_5_lutff_6_out_68600 = net_68600;
  assign seg_18_5_lutff_7_out_68601 = net_68601;
  assign seg_18_5_neigh_op_top_5_68722 = seg_18_6_lutff_5_out_68722;
  assign seg_18_5_neigh_op_top_6_68723 = seg_18_6_lutff_6_out_68723;
  assign seg_18_5_sp4_h_r_0_72560 = net_72560;
  assign seg_18_5_sp4_h_r_1_72561 = seg_21_5_sp4_h_r_36_72561;
  assign seg_18_5_sp4_h_r_2_72564 = net_72564;
  assign seg_18_5_sp4_h_r_4_72566 = seg_20_5_sp4_h_r_28_72566;
  assign seg_18_5_sp4_h_r_5_72567 = seg_21_5_sp4_h_r_40_72567;
  assign seg_18_5_sp4_h_r_9_72571 = seg_21_5_sp4_h_r_44_72571;
  assign seg_18_5_sp4_v_b_20_68503 = seg_18_3_sp4_v_b_44_68503;
  assign seg_18_6_lutff_1_out_68718 = net_68718;
  assign seg_18_6_lutff_3_out_68720 = net_68720;
  assign seg_18_6_lutff_5_out_68722 = net_68722;
  assign seg_18_6_lutff_6_out_68723 = net_68723;
  assign seg_18_6_lutff_7_out_68724 = net_68724;
  assign seg_18_6_neigh_op_bnl_5_64768 = seg_17_5_lutff_5_out_64768;
  assign seg_18_6_neigh_op_bot_2_68596 = seg_18_5_lutff_2_out_68596;
  assign seg_18_6_sp4_h_l_39_57364 = seg_14_6_sp4_h_r_2_57364;
  assign seg_18_6_sp4_h_l_45_57370 = seg_14_6_sp4_h_r_8_57370;
  assign seg_18_6_sp4_h_r_5_72690 = seg_21_6_sp4_h_r_40_72690;
  assign seg_18_6_sp4_h_r_7_72692 = seg_21_6_sp4_h_r_42_72692;
  assign seg_18_6_sp4_h_r_8_72693 = seg_20_6_sp4_h_r_32_72693;
  assign seg_18_6_sp4_r_v_b_15_72452 = net_72452;
  assign seg_18_6_sp4_v_b_0_68496 = net_68496;
  assign seg_18_6_sp4_v_b_8_68504 = net_68504;
  assign seg_18_7_neigh_op_bot_7_68724 = seg_18_6_lutff_7_out_68724;
  assign seg_18_7_sp12_h_r_14_45988 = net_45988;
  assign seg_18_7_sp12_h_r_16_42156 = net_42156;
  assign seg_18_7_sp12_h_r_18_38326 = net_38326;
  assign seg_18_7_sp12_v_b_18_72435 = net_72435;
  assign seg_18_7_sp4_h_l_43_57491 = seg_16_7_sp4_h_r_30_57491;
  assign seg_18_7_sp4_h_r_11_72809 = seg_21_7_sp4_h_r_46_72809;
  assign seg_18_7_sp4_h_r_14_68980 = net_68980;
  assign seg_18_7_sp4_h_r_20_68986 = net_68986;
  assign seg_18_7_sp4_h_r_28_65150 = net_65150;
  assign seg_18_7_sp4_h_r_2_72810 = net_72810;
  assign seg_18_7_sp4_h_r_3_72811 = seg_21_7_sp4_h_r_38_72811;
  assign seg_18_7_sp4_h_r_40_61320 = net_61320;
  assign seg_18_7_sp4_h_r_42_61322 = net_61322;
  assign seg_18_7_sp4_h_r_46_61316 = seg_16_7_sp4_h_r_22_61316;
  assign seg_18_7_sp4_r_v_b_10_72460 = seg_18_4_sp4_r_v_b_47_72460;
  assign seg_18_7_sp4_r_v_b_8_72458 = seg_18_4_sp4_r_v_b_45_72458;
  assign seg_18_7_sp4_v_b_14_68743 = net_68743;
  assign seg_18_7_sp4_v_b_1_68618 = seg_18_4_sp4_v_b_36_68618;
  assign seg_18_7_sp4_v_b_24_68865 = net_68865;
  assign seg_18_7_sp4_v_b_28_68869 = net_68869;
  assign seg_18_7_sp4_v_b_34_68875 = net_68875;
  assign seg_18_7_sp4_v_b_36_68987 = net_68987;
  assign seg_18_7_sp4_v_b_38_68989 = net_68989;
  assign seg_18_7_sp4_v_b_3_68620 = seg_18_4_sp4_v_b_38_68620;
  assign seg_18_7_sp4_v_b_42_68993 = net_68993;
  assign seg_18_7_sp4_v_b_44_68995 = net_68995;
  assign seg_18_7_sp4_v_b_46_68997 = seg_17_10_sp4_r_v_b_11_68997;
  assign seg_18_7_sp4_v_b_5_68622 = seg_18_4_sp4_v_b_40_68622;
  assign seg_18_7_sp4_v_b_7_68624 = seg_18_4_sp4_v_b_42_68624;
  assign seg_18_8_sp4_h_r_0_72929 = net_72929;
  assign seg_18_8_sp4_h_r_18_69107 = net_69107;
  assign seg_18_8_sp4_h_r_2_72933 = net_72933;
  assign seg_18_8_sp4_h_r_32_65277 = net_65277;
  assign seg_18_8_sp4_h_r_40_61443 = net_61443;
  assign seg_18_8_sp4_h_r_46_61439 = net_61439;
  assign seg_18_8_sp4_h_r_5_72936 = seg_21_8_sp4_h_r_40_72936;
  assign seg_18_8_sp4_h_r_9_72940 = seg_21_8_sp4_h_r_44_72940;
  assign seg_18_8_sp4_r_v_b_19_72702 = net_72702;
  assign seg_18_8_sp4_v_b_10_68752 = net_68752;
  assign seg_18_8_sp4_v_b_32_68996 = net_68996;
  assign seg_18_8_sp4_v_b_35_68997 = seg_17_10_sp4_r_v_b_11_68997;
  assign seg_18_8_sp4_v_b_3_68743 = seg_18_7_sp4_v_b_14_68743;
  assign seg_18_9_lutff_0_out_69086 = net_69086;
  assign seg_18_9_lutff_5_out_69091 = net_69091;
  assign seg_18_9_lutff_6_out_69092 = net_69092;
  assign seg_18_9_neigh_op_tnl_2_65380 = seg_17_10_lutff_2_out_65380;
  assign seg_18_9_neigh_op_top_4_69213 = seg_18_10_lutff_4_out_69213;
  assign seg_18_9_sp4_h_r_34_65392 = net_65392;
  assign seg_18_9_sp4_r_v_b_23_72829 = net_72829;
  assign seg_18_9_sp4_v_b_0_68865 = seg_18_7_sp4_v_b_24_68865;
  assign seg_18_9_sp4_v_b_10_68875 = seg_18_7_sp4_v_b_34_68875;
  assign seg_18_9_sp4_v_b_4_68869 = seg_18_7_sp4_v_b_28_68869;
  assign seg_19_0_span4_horz_r_12_64262 = net_64262;
  assign seg_19_0_span4_vert_12_72048 = net_72048;
  assign seg_19_10_sp4_v_b_10_72829 = seg_18_9_sp4_r_v_b_23_72829;
  assign seg_19_10_sp4_v_t_46_73320 = seg_18_14_sp4_r_v_b_11_73320;
  assign seg_19_11_sp4_v_b_8_72950 = seg_18_10_sp4_r_v_b_21_72950;
  assign seg_19_12_sp4_h_l_36_61929 = seg_16_12_sp4_h_r_12_61929;
  assign seg_19_17_sp4_h_l_38_62548 = seg_16_17_sp4_h_r_14_62548;
  assign seg_19_2_sp4_v_b_1_72048 = seg_19_0_span4_vert_12_72048;
  assign seg_19_4_sp4_h_l_43_60952 = seg_15_4_sp4_h_r_6_60952;
  assign seg_19_5_sp4_h_r_3_76290 = seg_22_5_sp4_h_r_38_76290;
  assign seg_19_5_sp4_h_r_5_76292 = seg_20_5_sp4_h_r_16_76292;
  assign seg_19_7_sp4_v_b_2_72452 = seg_18_6_sp4_r_v_b_15_72452;
  assign seg_19_8_sp4_h_r_1_76592 = seg_20_8_sp4_h_r_12_76592;
  assign seg_19_9_sp4_v_b_6_72702 = seg_18_8_sp4_r_v_b_19_72702;
  assign seg_1_10_lutff_0_out_1965 = net_1965;
  assign seg_1_10_lutff_1_out_1966 = net_1966;
  assign seg_1_10_lutff_3_out_1968 = net_1968;
  assign seg_1_10_lutff_4_out_1969 = net_1969;
  assign seg_1_10_lutff_5_out_1970 = net_1970;
  assign seg_1_10_lutff_6_out_1971 = net_1971;
  assign seg_1_10_lutff_7_out_1972 = net_1972;
  assign seg_1_10_neigh_op_tnr_1_8185 = seg_2_11_lutff_1_out_8185;
  assign seg_1_10_neigh_op_tnr_2_8186 = seg_2_11_lutff_2_out_8186;
  assign seg_1_10_neigh_op_tnr_6_8190 = seg_2_11_lutff_6_out_8190;
  assign seg_1_10_sp4_h_l_40_2273 = seg_0_10_sp4_h_r_40_2273;
  assign seg_1_10_sp4_h_r_12_2239 = net_2239;
  assign seg_1_10_sp4_h_r_4_8202 = net_8202;
  assign seg_1_10_sp4_r_v_b_13_7915 = net_7915;
  assign seg_1_10_sp4_r_v_b_29_8065 = net_8065;
  assign seg_1_10_sp4_r_v_b_5_7771 = net_7771;
  assign seg_1_10_sp4_v_b_6_1647 = seg_1_8_sp4_v_b_30_1647;
  assign seg_1_10_sp4_v_t_36_2492 = seg_0_12_sp4_r_v_b_25_2492;
  assign seg_1_10_sp4_v_t_42_2498 = seg_0_12_sp4_r_v_b_31_2498;
  assign seg_1_10_sp4_v_t_45_2501 = seg_0_13_sp4_r_v_b_21_2501;
  assign seg_1_11_lutff_0_out_2190 = net_2190;
  assign seg_1_11_lutff_1_out_2191 = net_2191;
  assign seg_1_11_lutff_2_out_2192 = net_2192;
  assign seg_1_11_lutff_4_out_2194 = net_2194;
  assign seg_1_11_lutff_5_out_2195 = net_2195;
  assign seg_1_11_lutff_7_out_2197 = net_2197;
  assign seg_1_11_neigh_op_rgt_3_8187 = seg_2_11_lutff_3_out_8187;
  assign seg_1_11_sp4_h_l_46_2485 = seg_0_11_sp4_h_r_46_2485;
  assign seg_1_11_sp4_h_r_6_8351 = net_8351;
  assign seg_1_11_sp4_h_r_9_8354 = seg_4_11_sp4_h_r_44_8354;
  assign seg_1_11_sp4_r_v_b_23_8072 = net_8072;
  assign seg_1_11_sp4_r_v_b_7_7920 = net_7920;
  assign seg_1_11_sp4_v_b_10_1860 = seg_1_9_sp4_v_b_34_1860;
  assign seg_1_11_sp4_v_b_28_2291 = net_2291;
  assign seg_1_11_sp4_v_b_37_2493 = seg_1_14_sp4_v_b_0_2493;
  assign seg_1_11_sp4_v_b_3_1851 = seg_1_8_sp4_v_b_38_1851;
  assign seg_1_11_sp4_v_b_47_2503 = seg_1_14_sp4_v_b_10_2503;
  assign seg_1_11_sp4_v_b_5_1853 = seg_1_8_sp4_v_b_40_1853;
  assign seg_1_11_sp4_v_b_6_1856 = net_1856;
  assign seg_1_11_sp4_v_t_38_2702 = seg_0_13_sp4_r_v_b_27_2702;
  assign seg_1_11_sp4_v_t_39_2703 = seg_0_12_sp4_r_v_b_39_2703;
  assign seg_1_12_lutff_3_out_2399 = net_2399;
  assign seg_1_12_lutff_5_out_2401 = net_2401;
  assign seg_1_12_lutff_6_out_2402 = net_2402;
  assign seg_1_12_sp4_h_r_24_2657 = net_2657;
  assign seg_1_12_sp4_h_r_36_2670 = net_2670;
  assign seg_1_12_sp4_r_v_b_31_8361 = net_8361;
  assign seg_1_12_sp4_r_v_b_33_8363 = net_8363;
  assign seg_1_12_sp4_v_b_1_2076 = seg_1_9_sp4_v_b_36_2076;
  assign seg_1_12_sp4_v_b_28_2497 = seg_1_14_sp4_v_b_4_2497;
  assign seg_1_12_sp4_v_b_3_2078 = seg_1_9_sp4_v_b_38_2078;
  assign seg_1_12_sp4_v_t_40_2913 = seg_0_16_sp4_r_v_b_5_2913;
  assign seg_1_13_sp4_h_l_38_2893 = seg_0_13_sp4_h_r_38_2893;
  assign seg_1_13_sp4_h_r_0_8637 = net_8637;
  assign seg_1_13_sp4_h_r_22_2864 = net_2864;
  assign seg_1_13_sp4_h_r_26_2868 = net_2868;
  assign seg_1_13_sp4_h_r_28_2870 = net_2870;
  assign seg_1_13_sp4_h_r_2_8641 = net_8641;
  assign seg_1_13_sp4_h_r_30_2872 = net_2872;
  assign seg_1_13_sp4_h_r_4_8643 = net_8643;
  assign seg_1_13_sp4_h_r_8_8647 = net_8647;
  assign seg_1_13_sp4_v_b_0_2287 = seg_0_10_sp4_r_v_b_37_2287;
  assign seg_1_13_sp4_v_b_10_2297 = seg_0_10_sp4_r_v_b_47_2297;
  assign seg_1_13_sp4_v_b_2_2289 = seg_0_10_sp4_r_v_b_39_2289;
  assign seg_1_13_sp4_v_b_4_2291 = seg_1_11_sp4_v_b_28_2291;
  assign seg_1_13_sp4_v_b_6_2293 = seg_0_10_sp4_r_v_b_43_2293;
  assign seg_1_13_sp4_v_b_8_2295 = seg_0_10_sp4_r_v_b_45_2295;
  assign seg_1_13_sp4_v_t_39_3139 = seg_0_16_sp4_r_v_b_15_3139;
  assign seg_1_14_lutff_1_out_2814 = net_2814;
  assign seg_1_14_lutff_3_out_2816 = net_2816;
  assign seg_1_14_lutff_4_out_2817 = net_2817;
  assign seg_1_14_lutff_6_out_2819 = net_2819;
  assign seg_1_14_neigh_op_top_3_3028 = seg_1_15_lutff_3_out_3028;
  assign seg_1_14_neigh_op_top_5_3030 = seg_1_15_lutff_5_out_3030;
  assign seg_1_14_neigh_op_top_7_3032 = seg_1_15_lutff_7_out_3032;
  assign seg_1_14_sp4_r_v_b_15_8505 = net_8505;
  assign seg_1_14_sp4_v_b_0_2493 = net_2493;
  assign seg_1_14_sp4_v_b_10_2503 = net_2503;
  assign seg_1_14_sp4_v_b_4_2497 = net_2497;
  assign seg_1_14_sp4_v_t_38_3348 = seg_1_17_sp4_v_b_14_3348;
  assign seg_1_15_lutff_0_out_3025 = net_3025;
  assign seg_1_15_lutff_1_out_3026 = net_3026;
  assign seg_1_15_lutff_2_out_3027 = net_3027;
  assign seg_1_15_lutff_3_out_3028 = net_3028;
  assign seg_1_15_lutff_4_out_3029 = net_3029;
  assign seg_1_15_lutff_5_out_3030 = net_3030;
  assign seg_1_15_lutff_6_out_3031 = net_3031;
  assign seg_1_15_lutff_7_out_3032 = net_3032;
  assign seg_1_15_sp4_v_b_24_3137 = seg_0_16_sp4_r_v_b_13_3137;
  assign seg_1_15_sp4_v_b_41_3351 = seg_0_17_sp4_r_v_b_17_3351;
  assign seg_1_15_sp4_v_b_46_3356 = seg_0_18_sp4_r_v_b_11_3356;
  assign seg_1_15_sp4_v_t_40_3556 = seg_0_17_sp4_r_v_b_29_3556;
  assign seg_1_15_sp4_v_t_43_3559 = seg_0_18_sp4_r_v_b_19_3559;
  assign seg_1_15_sp4_v_t_46_3562 = seg_0_17_sp4_r_v_b_35_3562;
  assign seg_1_16_lutff_0_out_3250 = net_3250;
  assign seg_1_16_lutff_2_out_3252 = net_3252;
  assign seg_1_16_lutff_3_out_3253 = net_3253;
  assign seg_1_16_lutff_4_out_3254 = net_3254;
  assign seg_1_16_lutff_5_out_3255 = net_3255;
  assign seg_1_16_lutff_6_out_3256 = net_3256;
  assign seg_1_16_sp4_h_r_2_9082 = net_9082;
  assign seg_1_16_sp4_v_b_10_2920 = seg_0_15_sp4_r_v_b_23_2920;
  assign seg_1_16_sp4_v_b_29_3350 = seg_0_18_sp4_r_v_b_5_3350;
  assign seg_1_16_sp4_v_b_33_3354 = seg_0_18_sp4_r_v_b_9_3354;
  assign seg_1_16_sp4_v_b_37_3553 = seg_0_18_sp4_r_v_b_13_3553;
  assign seg_1_17_lutff_1_out_3457 = net_3457;
  assign seg_1_17_lutff_2_out_3458 = net_3458;
  assign seg_1_17_neigh_op_top_0_3664 = seg_1_18_lutff_0_out_3664;
  assign seg_1_17_neigh_op_top_1_3665 = seg_1_18_lutff_1_out_3665;
  assign seg_1_17_neigh_op_top_4_3668 = seg_1_18_lutff_4_out_3668;
  assign seg_1_17_sp12_v_b_1_7459 = seg_1_6_sp12_v_b_22_7459;
  assign seg_1_17_sp4_r_v_b_7_8802 = net_8802;
  assign seg_1_17_sp4_v_b_14_3348 = net_3348;
  assign seg_1_18_lutff_0_out_3664 = net_3664;
  assign seg_1_18_lutff_1_out_3665 = net_3665;
  assign seg_1_18_lutff_4_out_3668 = net_3668;
  assign seg_1_18_lutff_6_out_3670 = net_3670;
  assign seg_1_18_neigh_op_top_5_3878 = seg_1_19_lutff_5_out_3878;
  assign seg_1_18_neigh_op_top_7_3880 = seg_1_19_lutff_7_out_3880;
  assign seg_1_18_sp4_v_b_43_3976 = seg_1_21_sp4_v_b_6_3976;
  assign seg_1_19_lutff_0_out_3873 = net_3873;
  assign seg_1_19_lutff_5_out_3878 = net_3878;
  assign seg_1_19_lutff_7_out_3880 = net_3880;
  assign seg_1_19_neigh_op_top_1_4086 = seg_1_20_lutff_1_out_4086;
  assign seg_1_19_neigh_op_top_6_4091 = seg_1_20_lutff_6_out_4091;
  assign seg_1_19_neigh_op_top_7_4092 = seg_1_20_lutff_7_out_4092;
  assign seg_1_19_sp4_v_t_38_4425 = seg_0_23_sp4_r_v_b_3_4425;
  assign seg_1_19_sp4_v_t_40_4427 = seg_0_23_sp4_r_v_b_5_4427;
  assign seg_1_19_sp4_v_t_42_4429 = seg_0_23_sp4_r_v_b_7_4429;
  assign seg_1_19_sp4_v_t_44_4431 = seg_0_23_sp4_r_v_b_9_4431;
  assign seg_1_19_sp4_v_t_46_4433 = seg_0_23_sp4_r_v_b_11_4433;
  assign seg_1_1_lutff_2_out_103 = net_103;
  assign seg_1_1_lutff_5_out_106 = net_106;
  assign seg_1_1_lutff_6_out_107 = net_107;
  assign seg_1_1_lutff_7_out_108 = net_108;
  assign seg_1_1_neigh_op_top_3_119 = seg_1_2_lutff_3_out_119;
  assign seg_1_1_neigh_op_top_6_122 = seg_1_2_lutff_6_out_122;
  assign seg_1_1_sp4_h_r_20_250 = seg_3_1_sp4_h_r_44_250;
  assign seg_1_1_sp4_r_v_b_29_6871 = net_6871;
  assign seg_1_1_sp4_r_v_b_45_6889 = net_6889;
  assign seg_1_1_sp4_v_b_46_292 = net_292;
  assign seg_1_20_lutff_1_out_4086 = net_4086;
  assign seg_1_20_lutff_2_out_4087 = net_4087;
  assign seg_1_20_lutff_6_out_4091 = net_4091;
  assign seg_1_20_lutff_7_out_4092 = net_4092;
  assign seg_1_20_sp4_v_b_36_4423 = seg_1_22_sp4_v_b_12_4423;
  assign seg_1_20_sp4_v_t_36_4650 = seg_0_24_sp4_r_v_b_1_4650;
  assign seg_1_20_sp4_v_t_39_4653 = seg_0_23_sp4_r_v_b_15_4653;
  assign seg_1_20_sp4_v_t_40_4654 = seg_0_24_sp4_r_v_b_5_4654;
  assign seg_1_20_sp4_v_t_44_4658 = seg_0_24_sp4_r_v_b_9_4658;
  assign seg_1_20_sp4_v_t_46_4660 = seg_0_24_sp4_r_v_b_11_4660;
  assign seg_1_21_lutff_0_out_4312 = net_4312;
  assign seg_1_21_neigh_op_top_5_4544 = seg_1_22_lutff_5_out_4544;
  assign seg_1_21_sp4_v_b_6_3976 = net_3976;
  assign seg_1_21_sp4_v_t_38_4879 = seg_0_25_sp4_r_v_b_3_4879;
  assign seg_1_21_sp4_v_t_39_4880 = seg_0_24_sp4_r_v_b_15_4880;
  assign seg_1_21_sp4_v_t_40_4881 = seg_0_25_sp4_r_v_b_5_4881;
  assign seg_1_22_lutff_1_out_4540 = net_4540;
  assign seg_1_22_lutff_5_out_4544 = net_4544;
  assign seg_1_22_sp4_v_b_12_4423 = net_4423;
  assign seg_1_22_sp4_v_t_37_5088 = seg_0_25_sp4_r_v_b_13_5088;
  assign seg_1_22_sp4_v_t_40_5091 = seg_0_24_sp4_r_v_b_29_5091;
  assign seg_1_22_sp4_v_t_44_5095 = seg_0_26_sp4_r_v_b_9_5095;
  assign seg_1_22_sp4_v_t_46_5097 = seg_0_24_sp4_r_v_b_35_5097;
  assign seg_1_23_lutff_2_out_4768 = net_4768;
  assign seg_1_23_sp4_v_b_42_5093 = seg_0_26_sp4_r_v_b_7_5093;
  assign seg_1_23_sp4_v_t_41_5298 = seg_0_26_sp4_r_v_b_17_5298;
  assign seg_1_23_sp4_v_t_42_5299 = seg_0_25_sp4_r_v_b_31_5299;
  assign seg_1_23_sp4_v_t_45_5302 = seg_0_26_sp4_r_v_b_21_5302;
  assign seg_1_24_sp4_v_t_46_5511 = seg_0_26_sp4_r_v_b_35_5511;
  assign seg_1_2_lutff_1_out_117 = net_117;
  assign seg_1_2_lutff_2_out_118 = net_118;
  assign seg_1_2_lutff_3_out_119 = net_119;
  assign seg_1_2_lutff_4_out_120 = net_120;
  assign seg_1_2_lutff_5_out_121 = net_121;
  assign seg_1_2_lutff_6_out_122 = net_122;
  assign seg_1_2_lutff_7_out_123 = net_123;
  assign seg_1_2_neigh_op_bot_2_103 = seg_1_1_lutff_2_out_103;
  assign seg_1_2_neigh_op_bot_5_106 = seg_1_1_lutff_5_out_106;
  assign seg_1_2_neigh_op_rgt_1_6826 = seg_2_2_lutff_1_out_6826;
  assign seg_1_2_neigh_op_rgt_6_6831 = seg_2_2_lutff_6_out_6831;
  assign seg_1_2_neigh_op_rgt_7_6832 = seg_2_2_lutff_7_out_6832;
  assign seg_1_2_neigh_op_top_2_453 = seg_1_3_lutff_2_out_453;
  assign seg_1_2_neigh_op_top_5_456 = seg_1_3_lutff_5_out_456;
  assign seg_1_2_neigh_op_top_7_458 = seg_1_3_lutff_7_out_458;
  assign seg_1_2_sp4_h_r_28_523 = net_523;
  assign seg_1_2_sp4_r_v_b_31_6886 = seg_2_1_sp4_v_b_42_6886;
  assign seg_1_3_lutff_0_out_451 = net_451;
  assign seg_1_3_lutff_1_out_452 = net_452;
  assign seg_1_3_lutff_2_out_453 = net_453;
  assign seg_1_3_lutff_3_out_454 = net_454;
  assign seg_1_3_lutff_4_out_455 = net_455;
  assign seg_1_3_lutff_5_out_456 = net_456;
  assign seg_1_3_lutff_6_out_457 = net_457;
  assign seg_1_3_lutff_7_out_458 = net_458;
  assign seg_1_3_neigh_op_bnr_0_6825 = seg_2_2_lutff_0_out_6825;
  assign seg_1_3_neigh_op_bot_5_121 = seg_1_2_lutff_5_out_121;
  assign seg_1_3_neigh_op_tnr_1_7156 = seg_2_4_lutff_1_out_7156;
  assign seg_1_3_neigh_op_top_1_679 = seg_1_4_lutff_1_out_679;
  assign seg_1_3_neigh_op_top_3_681 = seg_1_4_lutff_3_out_681;
  assign seg_1_3_sp4_h_r_10_7169 = net_7169;
  assign seg_1_3_sp4_h_r_20_788 = net_788;
  assign seg_1_3_sp4_h_r_38_761 = net_761;
  assign seg_1_3_sp4_h_r_8_7177 = net_7177;
  assign seg_1_3_sp4_r_v_b_21_6889 = seg_1_1_sp4_r_v_b_45_6889;
  assign seg_1_4_lutff_1_out_679 = net_679;
  assign seg_1_4_lutff_2_out_680 = net_680;
  assign seg_1_4_lutff_3_out_681 = net_681;
  assign seg_1_4_lutff_4_out_682 = net_682;
  assign seg_1_4_lutff_5_out_683 = net_683;
  assign seg_1_4_lutff_6_out_684 = net_684;
  assign seg_1_4_lutff_7_out_685 = net_685;
  assign seg_1_4_neigh_op_bot_0_451 = seg_1_3_lutff_0_out_451;
  assign seg_1_4_neigh_op_bot_1_452 = seg_1_3_lutff_1_out_452;
  assign seg_1_4_neigh_op_bot_3_454 = seg_1_3_lutff_3_out_454;
  assign seg_1_4_neigh_op_rgt_1_7156 = seg_2_4_lutff_1_out_7156;
  assign seg_1_4_neigh_op_rgt_2_7157 = seg_2_4_lutff_2_out_7157;
  assign seg_1_4_neigh_op_rgt_6_7161 = seg_2_4_lutff_6_out_7161;
  assign seg_1_4_neigh_op_tnr_2_7304 = seg_2_5_lutff_2_out_7304;
  assign seg_1_4_neigh_op_top_5_910 = seg_1_5_lutff_5_out_910;
  assign seg_1_4_sp4_v_b_11_292 = seg_1_1_sp4_v_b_46_292;
  assign seg_1_4_sp4_v_t_37_1227 = seg_0_7_sp4_r_v_b_13_1227;
  assign seg_1_5_lutff_0_out_905 = net_905;
  assign seg_1_5_lutff_5_out_910 = net_910;
  assign seg_1_5_lutff_6_out_911 = net_911;
  assign seg_1_5_neigh_op_bot_6_684 = seg_1_4_lutff_6_out_684;
  assign seg_1_5_neigh_op_rgt_4_7306 = seg_2_5_lutff_4_out_7306;
  assign seg_1_5_neigh_op_rgt_7_7309 = seg_2_5_lutff_7_out_7309;
  assign seg_1_5_sp4_h_l_38_1210 = seg_0_5_sp4_h_r_38_1210;
  assign seg_1_5_sp4_h_r_10_7463 = seg_3_5_sp4_h_r_34_7463;
  assign seg_1_5_sp4_h_r_14_1201 = net_1201;
  assign seg_1_5_sp4_h_r_18_1223 = net_1223;
  assign seg_1_5_sp4_h_r_20_1225 = net_1225;
  assign seg_1_5_sp4_h_r_22_1181 = net_1181;
  assign seg_1_5_sp4_h_r_6_7469 = seg_3_5_sp4_h_r_30_7469;
  assign seg_1_5_sp4_h_r_8_7471 = seg_3_5_sp4_h_r_32_7471;
  assign seg_1_5_sp4_r_v_b_1_7032 = net_7032;
  assign seg_1_5_sp4_v_b_24_1017 = net_1017;
  assign seg_1_5_sp4_v_b_34_1027 = net_1027;
  assign seg_1_5_sp4_v_b_42_1232 = seg_0_8_sp4_r_v_b_7_1232;
  assign seg_1_5_sp4_v_b_46_1236 = net_1236;
  assign seg_1_5_sp4_v_b_8_571 = net_571;
  assign seg_1_6_lutff_1_out_1131 = net_1131;
  assign seg_1_6_lutff_3_out_1133 = net_1133;
  assign seg_1_6_lutff_5_out_1135 = net_1135;
  assign seg_1_6_lutff_6_out_1136 = net_1136;
  assign seg_1_6_neigh_op_rgt_0_7449 = seg_2_6_lutff_0_out_7449;
  assign seg_1_6_neigh_op_rgt_3_7452 = seg_2_6_lutff_3_out_7452;
  assign seg_1_6_neigh_op_rgt_4_7453 = seg_2_6_lutff_4_out_7453;
  assign seg_1_6_sp12_v_b_22_7459 = net_7459;
  assign seg_1_6_sp4_h_l_44_1423 = seg_0_6_sp4_h_r_44_1423;
  assign seg_1_6_sp4_h_r_9_7619 = seg_2_6_sp4_h_r_20_7619;
  assign seg_1_6_sp4_v_b_40_1436 = net_1436;
  assign seg_1_6_sp4_v_b_44_1440 = net_1440;
  assign seg_1_6_sp4_v_b_8_798 = seg_0_5_sp4_r_v_b_21_798;
  assign seg_1_6_sp4_v_t_41_1645 = seg_0_7_sp4_r_v_b_41_1645;
  assign seg_1_7_lutff_1_out_1337 = net_1337;
  assign seg_1_7_sp4_h_r_2_7759 = seg_3_7_sp4_h_r_26_7759;
  assign seg_1_7_sp4_v_b_0_1017 = seg_1_5_sp4_v_b_24_1017;
  assign seg_1_7_sp4_v_b_10_1027 = seg_1_5_sp4_v_b_34_1027;
  assign seg_1_7_sp4_v_b_2_1019 = seg_0_6_sp4_r_v_b_15_1019;
  assign seg_1_7_sp4_v_b_6_1023 = seg_0_6_sp4_r_v_b_19_1023;
  assign seg_1_7_sp4_v_t_43_1856 = seg_1_11_sp4_v_b_6_1856;
  assign seg_1_8_lutff_0_out_1544 = net_1544;
  assign seg_1_8_lutff_1_out_1545 = net_1545;
  assign seg_1_8_lutff_2_out_1546 = net_1546;
  assign seg_1_8_lutff_3_out_1547 = net_1547;
  assign seg_1_8_lutff_4_out_1548 = net_1548;
  assign seg_1_8_lutff_6_out_1550 = net_1550;
  assign seg_1_8_lutff_7_out_1551 = net_1551;
  assign seg_1_8_sp12_h_r_0_7898 = seg_11_8_sp12_h_r_20_7898;
  assign seg_1_8_sp4_h_r_10_7904 = net_7904;
  assign seg_1_8_sp4_v_b_16_1436 = seg_1_6_sp4_v_b_40_1436;
  assign seg_1_8_sp4_v_b_30_1647 = net_1647;
  assign seg_1_8_sp4_v_b_38_1851 = net_1851;
  assign seg_1_8_sp4_v_b_3_1228 = seg_0_6_sp4_r_v_b_27_1228;
  assign seg_1_8_sp4_v_b_40_1853 = net_1853;
  assign seg_1_8_sp4_v_b_6_1233 = seg_0_7_sp4_r_v_b_19_1233;
  assign seg_1_8_sp4_v_b_8_1235 = seg_0_7_sp4_r_v_b_21_1235;
  assign seg_1_8_sp4_v_t_46_2086 = seg_0_12_sp4_r_v_b_11_2086;
  assign seg_1_9_lutff_5_out_1758 = net_1758;
  assign seg_1_9_lutff_7_out_1760 = net_1760;
  assign seg_1_9_neigh_op_top_0_1965 = seg_1_10_lutff_0_out_1965;
  assign seg_1_9_sp12_h_r_13_1992 = seg_6_9_sp12_h_r_22_1992;
  assign seg_1_9_sp12_h_r_5_2002 = seg_6_9_sp12_h_r_14_2002;
  assign seg_1_9_sp4_h_r_16_2071 = net_2071;
  assign seg_1_9_sp4_r_v_b_29_7918 = net_7918;
  assign seg_1_9_sp4_r_v_b_41_8066 = net_8066;
  assign seg_1_9_sp4_r_v_b_45_8070 = net_8070;
  assign seg_1_9_sp4_v_b_24_1850 = net_1850;
  assign seg_1_9_sp4_v_b_32_1858 = net_1858;
  assign seg_1_9_sp4_v_b_34_1860 = net_1860;
  assign seg_1_9_sp4_v_b_36_2076 = net_2076;
  assign seg_1_9_sp4_v_b_38_2078 = net_2078;
  assign seg_1_9_sp4_v_b_9_1440 = seg_1_6_sp4_v_b_44_1440;
  assign seg_1_9_sp4_v_t_38_2288 = seg_0_13_sp4_r_v_b_3_2288;
  assign seg_1_9_sp4_v_t_41_2291 = seg_1_11_sp4_v_b_28_2291;
  assign seg_20_10_lutff_0_out_76651 = net_76651;
  assign seg_20_10_lutff_1_out_76652 = net_76652;
  assign seg_20_10_lutff_5_out_76656 = net_76656;
  assign seg_20_10_neigh_op_bot_7_76556 = seg_20_9_lutff_7_out_76556;
  assign seg_20_10_neigh_op_top_6_76759 = seg_20_11_lutff_6_out_76759;
  assign seg_20_10_sp4_h_l_39_65517 = seg_18_10_sp4_h_r_26_65517;
  assign seg_20_10_sp4_h_l_43_65521 = seg_18_10_sp4_h_r_30_65521;
  assign seg_20_10_sp4_h_r_24_73175 = net_73175;
  assign seg_20_10_sp4_h_r_26_73179 = net_73179;
  assign seg_20_10_sp4_h_r_8_80216 = seg_22_10_sp4_h_r_32_80216;
  assign seg_20_10_sp4_v_b_11_76511 = seg_20_9_sp4_v_b_22_76511;
  assign seg_20_11_lutff_6_out_76759 = net_76759;
  assign seg_20_11_neigh_op_bot_1_76652 = seg_20_10_lutff_1_out_76652;
  assign seg_20_11_sp4_h_r_30_73306 = net_73306;
  assign seg_20_12_sp4_v_b_4_76710 = net_76710;
  assign seg_20_14_sp4_h_r_38_69841 = net_69841;
  assign seg_20_2_lutff_2_out_75801 = net_75801;
  assign seg_20_2_lutff_7_out_75806 = net_75806;
  assign seg_20_2_sp4_h_l_38_64534 = seg_17_2_sp4_h_r_14_64534;
  assign seg_20_2_sp4_h_r_36_68361 = net_68361;
  assign seg_20_2_sp4_h_r_46_68363 = net_68363;
  assign seg_20_3_lutff_0_out_75937 = net_75937;
  assign seg_20_3_lutff_1_out_75938 = net_75938;
  assign seg_20_3_neigh_op_rgt_3_79213 = seg_21_3_lutff_3_out_79213;
  assign seg_20_3_sp4_h_l_41_64658 = seg_16_3_sp4_h_r_4_64658;
  assign seg_20_3_sp4_h_l_43_64660 = seg_16_3_sp4_h_r_6_64660;
  assign seg_20_3_sp4_h_r_28_72320 = net_72320;
  assign seg_20_3_sp4_h_r_38_68488 = net_68488;
  assign seg_20_3_sp4_h_r_42_68492 = net_68492;
  assign seg_20_3_sp4_h_r_46_68486 = net_68486;
  assign seg_20_4_sp4_h_r_18_76192 = net_76192;
  assign seg_20_4_sp4_h_r_5_79475 = seg_21_4_sp4_h_r_16_79475;
  assign seg_20_4_sp4_h_r_7_79477 = seg_21_4_sp4_h_r_18_79477;
  assign seg_20_4_sp4_r_v_b_19_79241 = net_79241;
  assign seg_20_5_sp4_h_r_16_76292 = net_76292;
  assign seg_20_5_sp4_h_r_28_72566 = net_72566;
  assign seg_20_5_sp4_h_r_2_79595 = net_79595;
  assign seg_20_5_sp4_h_r_36_68730 = net_68730;
  assign seg_20_5_sp4_h_r_38_68734 = net_68734;
  assign seg_20_5_sp4_h_r_40_68736 = net_68736;
  assign seg_20_5_sp4_h_r_42_68738 = net_68738;
  assign seg_20_5_sp4_h_r_46_68732 = net_68732;
  assign seg_20_5_sp4_h_r_5_79598 = seg_23_5_sp4_h_r_40_79598;
  assign seg_20_5_sp4_h_r_8_79601 = seg_22_5_sp4_h_r_32_79601;
  assign seg_20_6_sp4_h_r_32_72693 = net_72693;
  assign seg_20_6_sp4_h_r_3_79719 = seg_21_6_sp4_h_r_14_79719;
  assign seg_20_6_sp4_h_r_40_68859 = net_68859;
  assign seg_20_6_sp4_v_b_26_76300 = net_76300;
  assign seg_20_6_sp4_v_t_41_76506 = seg_20_8_sp4_v_b_28_76506;
  assign seg_20_7_sp4_h_r_42_68984 = net_68984;
  assign seg_20_8_neigh_op_tnr_3_79951 = seg_21_9_lutff_3_out_79951;
  assign seg_20_8_sp4_h_r_12_76592 = net_76592;
  assign seg_20_8_sp4_v_b_28_76506 = net_76506;
  assign seg_20_8_sp4_v_b_2_76300 = seg_20_6_sp4_v_b_26_76300;
  assign seg_20_8_sp4_v_t_41_76710 = seg_20_12_sp4_v_b_4_76710;
  assign seg_20_9_lutff_7_out_76556 = net_76556;
  assign seg_20_9_neigh_op_bnr_1_79826 = seg_21_8_lutff_1_out_79826;
  assign seg_20_9_neigh_op_bnr_7_79832 = seg_21_8_lutff_7_out_79832;
  assign seg_20_9_neigh_op_rgt_7_79955 = seg_21_9_lutff_7_out_79955;
  assign seg_20_9_sp4_h_l_47_65392 = seg_18_9_sp4_h_r_34_65392;
  assign seg_20_9_sp4_h_r_42_69230 = net_69230;
  assign seg_20_9_sp4_h_r_8_80093 = net_80093;
  assign seg_20_9_sp4_h_r_9_80094 = seg_21_9_sp4_h_r_20_80094;
  assign seg_20_9_sp4_v_b_22_76511 = net_76511;
  assign seg_21_10_lutff_2_out_80073 = net_80073;
  assign seg_21_10_lutff_3_out_80074 = net_80074;
  assign seg_21_10_neigh_op_bot_0_79948 = seg_21_9_lutff_0_out_79948;
  assign seg_21_10_neigh_op_lft_0_76651 = seg_20_10_lutff_0_out_76651;
  assign seg_21_10_neigh_op_lft_5_76656 = seg_20_10_lutff_5_out_76656;
  assign seg_21_10_sp4_h_r_0_84037 = net_84037;
  assign seg_21_10_sp4_h_r_2_84041 = net_84041;
  assign seg_21_10_sp4_h_r_40_73182 = net_73182;
  assign seg_21_10_sp4_v_b_2_79852 = seg_21_8_sp4_v_b_26_79852;
  assign seg_21_10_sp4_v_b_7_79855 = seg_21_9_sp4_v_b_18_79855;
  assign seg_21_2_sp4_h_l_37_68360 = seg_17_2_sp4_h_r_0_68360;
  assign seg_21_3_lutff_3_out_79213 = net_79213;
  assign seg_21_3_neigh_op_rgt_0_83041 = seg_22_3_lutff_0_out_83041;
  assign seg_21_3_neigh_op_rgt_2_83043 = seg_22_3_lutff_2_out_83043;
  assign seg_21_3_neigh_op_tnr_6_83170 = seg_22_4_lutff_6_out_83170;
  assign seg_21_3_sp4_h_r_0_83176 = net_83176;
  assign seg_21_3_sp4_h_r_36_72315 = net_72315;
  assign seg_21_3_sp4_h_r_46_72317 = net_72317;
  assign seg_21_4_neigh_op_rgt_7_83171 = seg_22_4_lutff_7_out_83171;
  assign seg_21_4_neigh_op_tnr_6_83293 = seg_22_5_lutff_6_out_83293;
  assign seg_21_4_sp4_h_r_16_79475 = net_79475;
  assign seg_21_4_sp4_h_r_18_79477 = net_79477;
  assign seg_21_4_sp4_h_r_36_72438 = net_72438;
  assign seg_21_4_sp4_h_r_42_72446 = net_72446;
  assign seg_21_4_sp4_h_r_46_72440 = net_72440;
  assign seg_21_5_neigh_op_rgt_4_83291 = seg_22_5_lutff_4_out_83291;
  assign seg_21_5_sp4_h_r_36_72561 = net_72561;
  assign seg_21_5_sp4_h_r_3_83427 = seg_22_5_sp4_h_r_14_83427;
  assign seg_21_5_sp4_h_r_40_72567 = net_72567;
  assign seg_21_5_sp4_h_r_44_72571 = net_72571;
  assign seg_21_5_sp4_v_b_6_79241 = seg_20_4_sp4_r_v_b_19_79241;
  assign seg_21_6_lutff_6_out_79585 = net_79585;
  assign seg_21_6_neigh_op_rgt_4_83414 = seg_22_6_lutff_4_out_83414;
  assign seg_21_6_sp4_h_r_14_79719 = net_79719;
  assign seg_21_6_sp4_h_r_1_83546 = seg_22_6_sp4_h_r_12_83546;
  assign seg_21_6_sp4_h_r_40_72690 = net_72690;
  assign seg_21_6_sp4_h_r_42_72692 = net_72692;
  assign seg_21_7_lutff_1_out_79703 = net_79703;
  assign seg_21_7_lutff_2_out_79704 = net_79704;
  assign seg_21_7_neigh_op_tnr_2_83658 = seg_22_8_lutff_2_out_83658;
  assign seg_21_7_sp4_h_l_38_68980 = seg_18_7_sp4_h_r_14_68980;
  assign seg_21_7_sp4_h_r_38_72811 = net_72811;
  assign seg_21_7_sp4_h_r_46_72809 = net_72809;
  assign seg_21_8_lutff_1_out_79826 = net_79826;
  assign seg_21_8_lutff_7_out_79832 = net_79832;
  assign seg_21_8_neigh_op_bnr_2_83535 = seg_22_7_lutff_2_out_83535;
  assign seg_21_8_neigh_op_bnr_4_83537 = seg_22_7_lutff_4_out_83537;
  assign seg_21_8_neigh_op_bnr_5_83538 = seg_22_7_lutff_5_out_83538;
  assign seg_21_8_neigh_op_bnr_7_83540 = seg_22_7_lutff_7_out_83540;
  assign seg_21_8_neigh_op_bot_1_79703 = seg_21_7_lutff_1_out_79703;
  assign seg_21_8_neigh_op_bot_2_79704 = seg_21_7_lutff_2_out_79704;
  assign seg_21_8_neigh_op_rgt_0_83656 = seg_22_8_lutff_0_out_83656;
  assign seg_21_8_neigh_op_rgt_3_83659 = seg_22_8_lutff_3_out_83659;
  assign seg_21_8_neigh_op_rgt_4_83660 = seg_22_8_lutff_4_out_83660;
  assign seg_21_8_neigh_op_rgt_5_83661 = seg_22_8_lutff_5_out_83661;
  assign seg_21_8_neigh_op_rgt_6_83662 = seg_22_8_lutff_6_out_83662;
  assign seg_21_8_neigh_op_tnr_4_83783 = seg_22_9_lutff_4_out_83783;
  assign seg_21_8_neigh_op_tnr_6_83785 = seg_22_9_lutff_6_out_83785;
  assign seg_21_8_neigh_op_tnr_7_83786 = seg_22_9_lutff_7_out_83786;
  assign seg_21_8_neigh_op_top_6_79954 = seg_21_9_lutff_6_out_79954;
  assign seg_21_8_sp12_h_r_12_61432 = net_61432;
  assign seg_21_8_sp12_h_r_14_57603 = net_57603;
  assign seg_21_8_sp4_h_r_40_72936 = net_72936;
  assign seg_21_8_sp4_h_r_44_72940 = net_72940;
  assign seg_21_8_sp4_h_r_6_83799 = seg_23_8_sp4_h_r_30_83799;
  assign seg_21_8_sp4_v_b_26_79852 = net_79852;
  assign seg_21_9_lutff_0_out_79948 = net_79948;
  assign seg_21_9_lutff_3_out_79951 = net_79951;
  assign seg_21_9_lutff_4_out_79952 = net_79952;
  assign seg_21_9_lutff_6_out_79954 = net_79954;
  assign seg_21_9_lutff_7_out_79955 = net_79955;
  assign seg_21_9_neigh_op_bnr_5_83661 = seg_22_8_lutff_5_out_83661;
  assign seg_21_9_neigh_op_rgt_0_83779 = seg_22_9_lutff_0_out_83779;
  assign seg_21_9_neigh_op_rgt_3_83782 = seg_22_9_lutff_3_out_83782;
  assign seg_21_9_neigh_op_top_2_80073 = seg_21_10_lutff_2_out_80073;
  assign seg_21_9_neigh_op_top_3_80074 = seg_21_10_lutff_3_out_80074;
  assign seg_21_9_sp4_h_r_14_80088 = seg_23_9_sp4_h_r_38_80088;
  assign seg_21_9_sp4_h_r_20_80094 = net_80094;
  assign seg_21_9_sp4_v_b_18_79855 = net_79855;
  assign seg_22_10_sp12_h_r_18_54019 = seg_14_10_sp12_h_r_2_54019;
  assign seg_22_10_sp4_h_l_39_73179 = seg_20_10_sp4_h_r_26_73179;
  assign seg_22_10_sp4_h_r_11_87871 = seg_25_10_sp4_h_r_46_87871;
  assign seg_22_10_sp4_h_r_1_87869 = seg_25_10_sp4_h_r_36_87869;
  assign seg_22_10_sp4_h_r_32_80216 = net_80216;
  assign seg_22_10_sp4_h_r_3_87873 = seg_25_10_sp4_h_r_38_87873;
  assign seg_22_11_sp4_h_r_11_87994 = seg_25_11_sp4_h_r_46_87994;
  assign seg_22_11_sp4_h_r_1_87992 = seg_25_11_sp4_h_r_36_87992;
  assign seg_22_12_sp4_h_r_11_88117 = seg_25_12_sp4_h_r_46_88117;
  assign seg_22_12_sp4_h_r_5_88121 = seg_25_12_sp4_h_r_40_88121;
  assign seg_22_13_sp4_h_r_3_88242 = seg_25_13_sp4_h_r_38_88242;
  assign seg_22_13_sp4_h_r_5_88244 = seg_25_13_sp4_h_r_40_88244;
  assign seg_22_13_sp4_h_r_9_88248 = seg_25_13_sp4_h_r_44_88248;
  assign seg_22_3_lutff_0_out_83041 = net_83041;
  assign seg_22_3_lutff_2_out_83043 = net_83043;
  assign seg_22_3_sp4_h_r_8_87017 = net_87017;
  assign seg_22_4_lutff_6_out_83170 = net_83170;
  assign seg_22_4_lutff_7_out_83171 = net_83171;
  assign seg_22_4_neigh_op_tnr_7_87125 = seg_23_5_lutff_7_out_87125;
  assign seg_22_4_sp12_h_r_12_64771 = net_64771;
  assign seg_22_5_lutff_4_out_83291 = net_83291;
  assign seg_22_5_lutff_6_out_83293 = net_83293;
  assign seg_22_5_neigh_op_rgt_0_87118 = seg_23_5_lutff_0_out_87118;
  assign seg_22_5_neigh_op_rgt_1_87119 = seg_23_5_lutff_1_out_87119;
  assign seg_22_5_neigh_op_tnr_3_87244 = seg_23_6_lutff_3_out_87244;
  assign seg_22_5_sp4_h_r_11_87256 = seg_25_5_sp4_h_r_46_87256;
  assign seg_22_5_sp4_h_r_14_83427 = net_83427;
  assign seg_22_5_sp4_h_r_1_87254 = seg_25_5_sp4_h_r_36_87254;
  assign seg_22_5_sp4_h_r_32_79601 = net_79601;
  assign seg_22_5_sp4_h_r_38_76290 = net_76290;
  assign seg_22_5_sp4_h_r_3_87258 = seg_25_5_sp4_h_r_38_87258;
  assign seg_22_5_sp4_h_r_7_87262 = seg_25_5_sp4_h_r_42_87262;
  assign seg_22_5_sp4_h_r_9_87264 = seg_25_5_sp4_h_r_44_87264;
  assign seg_22_6_lutff_4_out_83414 = net_83414;
  assign seg_22_6_neigh_op_rgt_7_87248 = seg_23_6_lutff_7_out_87248;
  assign seg_22_6_sp12_h_r_16_57356 = seg_14_6_sp12_h_r_0_57356;
  assign seg_22_6_sp4_h_r_12_83546 = net_83546;
  assign seg_22_6_sp4_h_r_1_87377 = seg_25_6_sp4_h_r_36_87377;
  assign seg_22_6_sp4_h_r_5_87383 = seg_25_6_sp4_h_r_40_87383;
  assign seg_22_7_lutff_2_out_83535 = net_83535;
  assign seg_22_7_lutff_4_out_83537 = net_83537;
  assign seg_22_7_lutff_5_out_83538 = net_83538;
  assign seg_22_7_lutff_7_out_83540 = net_83540;
  assign seg_22_7_sp4_h_r_11_87502 = seg_25_7_sp4_h_r_46_87502;
  assign seg_22_7_sp4_h_r_7_87508 = seg_25_7_sp4_h_r_42_87508;
  assign seg_22_7_sp4_h_r_9_87510 = seg_25_7_sp4_h_r_44_87510;
  assign seg_22_8_lutff_0_out_83656 = net_83656;
  assign seg_22_8_lutff_2_out_83658 = net_83658;
  assign seg_22_8_lutff_3_out_83659 = net_83659;
  assign seg_22_8_lutff_4_out_83660 = net_83660;
  assign seg_22_8_lutff_5_out_83661 = net_83661;
  assign seg_22_8_lutff_6_out_83662 = net_83662;
  assign seg_22_8_sp4_h_r_5_87629 = seg_25_8_sp4_h_r_40_87629;
  assign seg_22_8_sp4_h_r_7_87631 = seg_25_8_sp4_h_r_42_87631;
  assign seg_22_8_sp4_h_r_9_87633 = seg_25_8_sp4_h_r_44_87633;
  assign seg_22_9_lutff_0_out_83779 = net_83779;
  assign seg_22_9_lutff_3_out_83782 = net_83782;
  assign seg_22_9_lutff_4_out_83783 = net_83783;
  assign seg_22_9_lutff_6_out_83785 = net_83785;
  assign seg_22_9_lutff_7_out_83786 = net_83786;
  assign seg_23_0_span4_vert_0_86737 = net_86737;
  assign seg_23_0_span4_vert_16_86745 = net_86745;
  assign seg_23_10_sp4_h_r_0_91699 = seg_25_10_sp4_h_r_24_91699;
  assign seg_23_10_sp4_h_r_10_91701 = seg_25_10_sp4_h_r_34_91701;
  assign seg_23_10_sp4_h_r_2_91703 = seg_25_10_sp4_h_r_26_91703;
  assign seg_23_10_sp4_h_r_4_91705 = seg_25_10_sp4_h_r_28_91705;
  assign seg_23_12_sp4_h_r_4_91951 = seg_25_12_sp4_h_r_28_91951;
  assign seg_23_13_sp4_h_r_6_92076 = seg_25_13_sp4_h_r_30_92076;
  assign seg_23_1_sp4_v_b_0_86737 = seg_23_0_span4_vert_0_86737;
  assign seg_23_2_sp4_v_b_5_86745 = seg_23_0_span4_vert_16_86745;
  assign seg_23_3_sp4_v_t_39_87145 = seg_23_5_sp4_v_b_26_87145;
  assign seg_23_4_sp4_h_l_42_76192 = seg_20_4_sp4_h_r_18_76192;
  assign seg_23_5_lutff_0_out_87118 = net_87118;
  assign seg_23_5_lutff_1_out_87119 = net_87119;
  assign seg_23_5_lutff_7_out_87125 = net_87125;
  assign seg_23_5_neigh_op_top_1_87242 = seg_23_6_lutff_1_out_87242;
  assign seg_23_5_sp4_h_r_0_91084 = seg_25_5_sp4_h_r_24_91084;
  assign seg_23_5_sp4_h_r_40_79598 = net_79598;
  assign seg_23_5_sp4_h_r_8_91094 = seg_25_5_sp4_h_r_32_91094;
  assign seg_23_5_sp4_v_b_26_87145 = net_87145;
  assign seg_23_6_lutff_1_out_87242 = net_87242;
  assign seg_23_6_lutff_3_out_87244 = net_87244;
  assign seg_23_6_lutff_7_out_87248 = net_87248;
  assign seg_23_6_sp4_h_r_10_91209 = seg_25_6_sp4_h_r_34_91209;
  assign seg_23_6_sp4_h_r_8_91217 = seg_25_6_sp4_h_r_32_91217;
  assign seg_23_7_sp4_h_r_0_91330 = seg_25_7_sp4_h_r_24_91330;
  assign seg_23_8_sp4_h_r_30_83799 = net_83799;
  assign seg_23_8_sp4_h_r_8_91463 = seg_25_8_sp4_h_r_32_91463;
  assign seg_23_9_sp4_h_r_38_80088 = net_80088;
  assign seg_24_13_sp4_h_r_9_96090 = seg_25_13_sp4_h_r_20_96090;
  assign seg_24_6_sp4_h_r_11_95109 = seg_25_6_sp4_h_r_22_95109;
  assign seg_24_6_sp4_h_r_1_95107 = seg_25_6_sp4_h_r_12_95107;
  assign seg_25_10_sp4_h_r_24_91699 = net_91699;
  assign seg_25_10_sp4_h_r_26_91703 = net_91703;
  assign seg_25_10_sp4_h_r_28_91705 = net_91705;
  assign seg_25_10_sp4_h_r_34_91701 = net_91701;
  assign seg_25_10_sp4_h_r_36_87869 = net_87869;
  assign seg_25_10_sp4_h_r_38_87873 = net_87873;
  assign seg_25_10_sp4_h_r_46_87871 = net_87871;
  assign seg_25_10_sp4_v_b_0_95258 = net_95258;
  assign seg_25_11_sp4_h_r_2_100240 = net_100240;
  assign seg_25_11_sp4_h_r_36_87992 = net_87992;
  assign seg_25_11_sp4_h_r_46_87994 = net_87994;
  assign seg_25_11_sp4_v_b_0_95397 = net_95397;
  assign seg_25_11_sp4_v_b_10_95407 = net_95407;
  assign seg_25_11_sp4_v_b_12_95535 = net_95535;
  assign seg_25_11_sp4_v_b_22_95545 = net_95545;
  assign seg_25_11_sp4_v_b_8_95405 = net_95405;
  assign seg_25_12_sp4_h_r_28_91951 = net_91951;
  assign seg_25_12_sp4_h_r_40_88121 = net_88121;
  assign seg_25_12_sp4_h_r_46_88117 = net_88117;
  assign seg_25_12_sp4_v_b_10_95546 = net_95546;
  assign seg_25_12_sp4_v_b_16_95678 = net_95678;
  assign seg_25_12_sp4_v_b_20_95682 = net_95682;
  assign seg_25_12_sp4_v_b_2_95538 = net_95538;
  assign seg_25_12_sp4_v_b_6_95542 = net_95542;
  assign seg_25_13_sp4_h_r_20_96090 = net_96090;
  assign seg_25_13_sp4_h_r_30_92076 = net_92076;
  assign seg_25_13_sp4_h_r_38_88242 = net_88242;
  assign seg_25_13_sp4_h_r_40_88244 = net_88244;
  assign seg_25_13_sp4_h_r_44_88248 = net_88248;
  assign seg_25_13_sp4_v_b_0_95675 = net_95675;
  assign seg_25_13_sp4_v_b_10_95685 = net_95685;
  assign seg_25_13_sp4_v_b_2_95677 = net_95677;
  assign seg_25_3_sp4_v_t_37_94841 = seg_25_7_sp4_v_b_0_94841;
  assign seg_25_3_sp4_v_t_39_94843 = seg_25_7_sp4_v_b_2_94843;
  assign seg_25_4_sp4_v_t_41_94984 = seg_25_8_sp4_v_b_4_94984;
  assign seg_25_4_sp4_v_t_43_94986 = seg_25_6_sp4_v_b_30_94986;
  assign seg_25_4_sp4_v_t_44_94987 = seg_25_7_sp4_v_b_20_94987;
  assign seg_25_5_sp4_h_r_24_91084 = net_91084;
  assign seg_25_5_sp4_h_r_32_91094 = net_91094;
  assign seg_25_5_sp4_h_r_36_87254 = net_87254;
  assign seg_25_5_sp4_h_r_38_87258 = net_87258;
  assign seg_25_5_sp4_h_r_42_87262 = net_87262;
  assign seg_25_5_sp4_h_r_44_87264 = net_87264;
  assign seg_25_5_sp4_h_r_46_87256 = net_87256;
  assign seg_25_5_sp4_v_b_34_94851 = net_94851;
  assign seg_25_5_sp4_v_t_42_95124 = seg_25_8_sp4_v_b_18_95124;
  assign seg_25_5_sp4_v_t_46_95128 = seg_25_8_sp4_v_b_22_95128;
  assign seg_25_6_sp4_h_r_10_99458 = net_99458;
  assign seg_25_6_sp4_h_r_12_95107 = net_95107;
  assign seg_25_6_sp4_h_r_22_95109 = net_95109;
  assign seg_25_6_sp4_h_r_32_91217 = net_91217;
  assign seg_25_6_sp4_h_r_34_91209 = net_91209;
  assign seg_25_6_sp4_h_r_36_87377 = net_87377;
  assign seg_25_6_sp4_h_r_40_87383 = net_87383;
  assign seg_25_6_sp4_v_b_30_94986 = net_94986;
  assign seg_25_6_sp4_v_t_38_95259 = seg_25_7_sp4_v_b_38_95259;
  assign seg_25_6_sp4_v_t_43_95264 = seg_25_8_sp4_v_b_30_95264;
  assign seg_25_7_sp4_h_r_24_91330 = net_91330;
  assign seg_25_7_sp4_h_r_42_87508 = net_87508;
  assign seg_25_7_sp4_h_r_44_87510 = net_87510;
  assign seg_25_7_sp4_h_r_46_87502 = net_87502;
  assign seg_25_7_sp4_v_b_0_94841 = net_94841;
  assign seg_25_7_sp4_v_b_10_94851 = seg_25_5_sp4_v_b_34_94851;
  assign seg_25_7_sp4_v_b_20_94987 = net_94987;
  assign seg_25_7_sp4_v_b_2_94843 = net_94843;
  assign seg_25_7_sp4_v_b_38_95259 = net_95259;
  assign seg_25_7_sp4_v_t_37_95397 = seg_25_11_sp4_v_b_0_95397;
  assign seg_25_7_sp4_v_t_45_95405 = seg_25_11_sp4_v_b_8_95405;
  assign seg_25_7_sp4_v_t_47_95407 = seg_25_11_sp4_v_b_10_95407;
  assign seg_25_8_sp4_h_r_32_91463 = net_91463;
  assign seg_25_8_sp4_h_r_40_87629 = net_87629;
  assign seg_25_8_sp4_h_r_42_87631 = net_87631;
  assign seg_25_8_sp4_h_r_44_87633 = net_87633;
  assign seg_25_8_sp4_v_b_18_95124 = net_95124;
  assign seg_25_8_sp4_v_b_22_95128 = net_95128;
  assign seg_25_8_sp4_v_b_30_95264 = net_95264;
  assign seg_25_8_sp4_v_b_4_94984 = net_94984;
  assign seg_25_8_sp4_v_t_36_95535 = seg_25_11_sp4_v_b_12_95535;
  assign seg_25_8_sp4_v_t_39_95538 = seg_25_12_sp4_v_b_2_95538;
  assign seg_25_8_sp4_v_t_43_95542 = seg_25_12_sp4_v_b_6_95542;
  assign seg_25_8_sp4_v_t_46_95545 = seg_25_11_sp4_v_b_22_95545;
  assign seg_25_8_sp4_v_t_47_95546 = seg_25_12_sp4_v_b_10_95546;
  assign seg_25_9_sp4_v_t_37_95675 = seg_25_13_sp4_v_b_0_95675;
  assign seg_25_9_sp4_v_t_39_95677 = seg_25_13_sp4_v_b_2_95677;
  assign seg_25_9_sp4_v_t_40_95678 = seg_25_12_sp4_v_b_16_95678;
  assign seg_25_9_sp4_v_t_44_95682 = seg_25_12_sp4_v_b_20_95682;
  assign seg_25_9_sp4_v_t_47_95685 = seg_25_13_sp4_v_b_10_95685;
  assign seg_2_10_lutff_0_out_8037 = net_8037;
  assign seg_2_10_lutff_2_out_8039 = net_8039;
  assign seg_2_10_lutff_4_out_8041 = net_8041;
  assign seg_2_10_lutff_6_out_8043 = net_8043;
  assign seg_2_10_lutff_7_out_8044 = net_8044;
  assign seg_2_10_neigh_op_lft_6_1971 = seg_1_10_lutff_6_out_1971;
  assign seg_2_10_neigh_op_tnl_0_2190 = seg_1_11_lutff_0_out_2190;
  assign seg_2_10_neigh_op_tnl_1_2191 = seg_1_11_lutff_1_out_2191;
  assign seg_2_10_neigh_op_tnl_4_2194 = seg_1_11_lutff_4_out_2194;
  assign seg_2_10_neigh_op_tnl_5_2195 = seg_1_11_lutff_5_out_2195;
  assign seg_2_10_sp4_h_r_2_12516 = seg_4_10_sp4_h_r_26_12516;
  assign seg_2_10_sp4_h_r_42_2248 = net_2248;
  assign seg_2_10_sp4_r_v_b_37_12525 = net_12525;
  assign seg_2_10_sp4_v_t_36_8355 = seg_2_13_sp4_v_b_12_8355;
  assign seg_2_10_sp4_v_t_42_8361 = seg_1_12_sp4_r_v_b_31_8361;
  assign seg_2_10_sp4_v_t_43_8362 = seg_2_14_sp4_v_b_6_8362;
  assign seg_2_10_sp4_v_t_44_8363 = seg_1_12_sp4_r_v_b_33_8363;
  assign seg_2_10_sp4_v_t_45_8364 = seg_2_14_sp4_v_b_8_8364;
  assign seg_2_11_lutff_1_out_8185 = net_8185;
  assign seg_2_11_lutff_2_out_8186 = net_8186;
  assign seg_2_11_lutff_3_out_8187 = net_8187;
  assign seg_2_11_lutff_5_out_8189 = net_8189;
  assign seg_2_11_lutff_6_out_8190 = net_8190;
  assign seg_2_11_neigh_op_bot_4_8041 = seg_2_10_lutff_4_out_8041;
  assign seg_2_11_neigh_op_tnr_1_12624 = seg_3_12_lutff_1_out_12624;
  assign seg_2_11_neigh_op_tnr_2_12625 = seg_3_12_lutff_2_out_12625;
  assign seg_2_11_neigh_op_tnr_3_12626 = seg_3_12_lutff_3_out_12626;
  assign seg_2_11_neigh_op_tnr_4_12627 = seg_3_12_lutff_4_out_12627;
  assign seg_2_11_neigh_op_tnr_5_12628 = seg_3_12_lutff_5_out_12628;
  assign seg_2_11_neigh_op_tnr_6_12629 = seg_3_12_lutff_6_out_12629;
  assign seg_2_11_neigh_op_tnr_7_12630 = seg_3_12_lutff_7_out_12630;
  assign seg_2_11_sp4_r_v_b_31_12530 = net_12530;
  assign seg_2_11_sp4_r_v_b_47_12658 = net_12658;
  assign seg_2_11_sp4_v_b_5_7918 = seg_1_9_sp4_r_v_b_29_7918;
  assign seg_2_11_sp4_v_b_8_7923 = net_7923;
  assign seg_2_11_sp4_v_t_39_8505 = seg_1_14_sp4_r_v_b_15_8505;
  assign seg_2_12_lutff_0_out_8331 = net_8331;
  assign seg_2_12_lutff_1_out_8332 = net_8332;
  assign seg_2_12_lutff_2_out_8333 = net_8333;
  assign seg_2_12_lutff_3_out_8334 = net_8334;
  assign seg_2_12_lutff_4_out_8335 = net_8335;
  assign seg_2_12_lutff_5_out_8336 = net_8336;
  assign seg_2_12_lutff_6_out_8337 = net_8337;
  assign seg_2_12_neigh_op_rgt_7_12630 = seg_3_12_lutff_7_out_12630;
  assign seg_2_12_sp4_h_l_36_2670 = seg_1_12_sp4_h_r_36_2670;
  assign seg_2_12_sp4_h_r_11_12761 = seg_5_12_sp4_h_r_46_12761;
  assign seg_2_12_sp4_r_v_b_31_12653 = net_12653;
  assign seg_2_12_sp4_v_b_10_8072 = seg_1_11_sp4_r_v_b_23_8072;
  assign seg_2_12_sp4_v_b_11_8071 = seg_2_9_sp4_v_b_46_8071;
  assign seg_2_12_sp4_v_b_4_8066 = seg_1_9_sp4_r_v_b_41_8066;
  assign seg_2_12_sp4_v_b_8_8070 = seg_1_9_sp4_r_v_b_45_8070;
  assign seg_2_13_lutff_0_out_8478 = net_8478;
  assign seg_2_13_lutff_1_out_8479 = net_8479;
  assign seg_2_13_lutff_4_out_8482 = net_8482;
  assign seg_2_13_lutff_6_out_8484 = net_8484;
  assign seg_2_13_lutff_7_out_8485 = net_8485;
  assign seg_2_13_neigh_op_bnr_7_12630 = seg_3_12_lutff_7_out_12630;
  assign seg_2_13_neigh_op_tnl_1_2814 = seg_1_14_lutff_1_out_2814;
  assign seg_2_13_neigh_op_tnl_3_2816 = seg_1_14_lutff_3_out_2816;
  assign seg_2_13_neigh_op_tnr_5_12874 = seg_3_14_lutff_5_out_12874;
  assign seg_2_13_sp4_h_l_37_2878 = seg_0_13_sp4_h_r_24_2878;
  assign seg_2_13_sp4_h_r_10_12883 = net_12883;
  assign seg_2_13_sp4_h_r_26_2873 = net_2873;
  assign seg_2_13_sp4_h_r_4_12887 = net_12887;
  assign seg_2_13_sp4_h_r_6_12889 = net_12889;
  assign seg_2_13_sp4_r_v_b_11_12534 = net_12534;
  assign seg_2_13_sp4_r_v_b_23_12658 = seg_2_11_sp4_r_v_b_47_12658;
  assign seg_2_13_sp4_v_b_10_8219 = net_8219;
  assign seg_2_13_sp4_v_b_12_8355 = net_8355;
  assign seg_2_13_sp4_v_t_42_8802 = seg_1_17_sp4_r_v_b_7_8802;
  assign seg_2_14_neigh_op_bnr_7_12753 = seg_3_13_lutff_7_out_12753;
  assign seg_2_14_neigh_op_rgt_0_12869 = seg_3_14_lutff_0_out_12869;
  assign seg_2_14_neigh_op_rgt_1_12870 = seg_3_14_lutff_1_out_12870;
  assign seg_2_14_neigh_op_top_1_8773 = seg_2_15_lutff_1_out_8773;
  assign seg_2_14_neigh_op_top_2_8774 = seg_2_15_lutff_2_out_8774;
  assign seg_2_14_neigh_op_top_3_8775 = seg_2_15_lutff_3_out_8775;
  assign seg_2_14_sp4_h_r_10_13006 = net_13006;
  assign seg_2_14_sp4_h_r_12_8785 = net_8785;
  assign seg_2_14_sp4_h_r_36_3092 = net_3092;
  assign seg_2_14_sp4_r_v_b_31_12899 = net_12899;
  assign seg_2_14_sp4_r_v_b_35_12903 = net_12903;
  assign seg_2_14_sp4_v_b_6_8362 = net_8362;
  assign seg_2_14_sp4_v_b_8_8364 = net_8364;
  assign seg_2_15_lutff_1_out_8773 = net_8773;
  assign seg_2_15_lutff_2_out_8774 = net_8774;
  assign seg_2_15_lutff_3_out_8775 = net_8775;
  assign seg_2_15_lutff_4_out_8776 = net_8776;
  assign seg_2_15_lutff_6_out_8778 = net_8778;
  assign seg_2_15_neigh_op_bnl_6_2819 = seg_1_14_lutff_6_out_2819;
  assign seg_2_15_neigh_op_lft_2_3027 = seg_1_15_lutff_2_out_3027;
  assign seg_2_15_neigh_op_tnl_3_3253 = seg_1_16_lutff_3_out_3253;
  assign seg_2_15_neigh_op_top_1_8920 = seg_2_16_lutff_1_out_8920;
  assign seg_2_15_neigh_op_top_2_8921 = seg_2_16_lutff_2_out_8921;
  assign seg_2_15_neigh_op_top_6_8925 = seg_2_16_lutff_6_out_8925;
  assign seg_2_15_neigh_op_top_7_8926 = seg_2_16_lutff_7_out_8926;
  assign seg_2_15_sp4_h_r_10_13129 = net_13129;
  assign seg_2_15_sp4_h_r_14_8936 = net_8936;
  assign seg_2_16_lutff_0_out_8919 = net_8919;
  assign seg_2_16_lutff_1_out_8920 = net_8920;
  assign seg_2_16_lutff_2_out_8921 = net_8921;
  assign seg_2_16_lutff_3_out_8922 = net_8922;
  assign seg_2_16_lutff_4_out_8923 = net_8923;
  assign seg_2_16_lutff_5_out_8924 = net_8924;
  assign seg_2_16_lutff_6_out_8925 = net_8925;
  assign seg_2_16_lutff_7_out_8926 = net_8926;
  assign seg_2_16_neigh_op_lft_2_3252 = seg_1_16_lutff_2_out_3252;
  assign seg_2_16_neigh_op_rgt_7_13122 = seg_3_16_lutff_7_out_13122;
  assign seg_2_16_neigh_op_tnl_1_3457 = seg_1_17_lutff_1_out_3457;
  assign seg_2_16_neigh_op_tnl_2_3458 = seg_1_17_lutff_2_out_3458;
  assign seg_2_16_neigh_op_top_2_9068 = seg_2_17_lutff_2_out_9068;
  assign seg_2_16_neigh_op_top_7_9073 = seg_2_17_lutff_7_out_9073;
  assign seg_2_16_sp4_v_b_43_9097 = seg_2_19_sp4_v_b_6_9097;
  assign seg_2_17_lutff_2_out_9068 = net_9068;
  assign seg_2_17_lutff_5_out_9071 = net_9071;
  assign seg_2_17_lutff_7_out_9073 = net_9073;
  assign seg_2_17_neigh_op_tnl_6_3670 = seg_1_18_lutff_6_out_3670;
  assign seg_2_17_neigh_op_top_4_9217 = seg_2_18_lutff_4_out_9217;
  assign seg_2_17_sp4_h_l_39_3731 = seg_0_17_sp4_h_r_26_3731;
  assign seg_2_17_sp4_v_t_39_9387 = seg_2_21_sp4_v_b_2_9387;
  assign seg_2_18_lutff_0_out_9213 = net_9213;
  assign seg_2_18_lutff_1_out_9214 = net_9214;
  assign seg_2_18_lutff_4_out_9217 = net_9217;
  assign seg_2_18_lutff_6_out_9219 = net_9219;
  assign seg_2_18_lutff_7_out_9220 = net_9220;
  assign seg_2_18_neigh_op_top_1_9361 = seg_2_19_lutff_1_out_9361;
  assign seg_2_18_neigh_op_top_5_9365 = seg_2_19_lutff_5_out_9365;
  assign seg_2_18_neigh_op_top_7_9367 = seg_2_19_lutff_7_out_9367;
  assign seg_2_19_lutff_0_out_9360 = net_9360;
  assign seg_2_19_lutff_1_out_9361 = net_9361;
  assign seg_2_19_lutff_4_out_9364 = net_9364;
  assign seg_2_19_lutff_5_out_9365 = net_9365;
  assign seg_2_19_lutff_6_out_9366 = net_9366;
  assign seg_2_19_lutff_7_out_9367 = net_9367;
  assign seg_2_19_neigh_op_lft_0_3873 = seg_1_19_lutff_0_out_3873;
  assign seg_2_19_neigh_op_top_3_9510 = seg_2_20_lutff_3_out_9510;
  assign seg_2_19_neigh_op_top_4_9511 = seg_2_20_lutff_4_out_9511;
  assign seg_2_19_neigh_op_top_5_9512 = seg_2_20_lutff_5_out_9512;
  assign seg_2_19_neigh_op_top_7_9514 = seg_2_20_lutff_7_out_9514;
  assign seg_2_19_sp4_v_b_6_9097 = net_9097;
  assign seg_2_1_lutff_0_out_6673 = net_6673;
  assign seg_2_1_lutff_1_out_6674 = net_6674;
  assign seg_2_1_lutff_3_out_6676 = net_6676;
  assign seg_2_1_lutff_5_out_6678 = net_6678;
  assign seg_2_1_lutff_7_out_6680 = net_6680;
  assign seg_2_1_neigh_op_rgt_6_11235 = seg_3_1_lutff_6_out_11235;
  assign seg_2_1_neigh_op_tnl_7_123 = seg_1_2_lutff_7_out_123;
  assign seg_2_1_neigh_op_top_4_6829 = seg_2_2_lutff_4_out_6829;
  assign seg_2_1_sp4_v_b_42_6886 = net_6886;
  assign seg_2_1_sp4_v_b_47_6891 = seg_2_4_sp4_v_b_10_6891;
  assign seg_2_20_lutff_1_out_9508 = net_9508;
  assign seg_2_20_lutff_3_out_9510 = net_9510;
  assign seg_2_20_lutff_4_out_9511 = net_9511;
  assign seg_2_20_lutff_5_out_9512 = net_9512;
  assign seg_2_20_lutff_7_out_9514 = net_9514;
  assign seg_2_20_neigh_op_lft_2_4087 = seg_1_20_lutff_2_out_4087;
  assign seg_2_20_neigh_op_tnl_0_4312 = seg_1_21_lutff_0_out_4312;
  assign seg_2_20_neigh_op_top_4_9658 = seg_2_21_lutff_4_out_9658;
  assign seg_2_21_lutff_4_out_9658 = net_9658;
  assign seg_2_21_neigh_op_top_0_9801 = seg_2_22_lutff_0_out_9801;
  assign seg_2_21_neigh_op_top_5_9806 = seg_2_22_lutff_5_out_9806;
  assign seg_2_21_sp4_v_b_2_9387 = net_9387;
  assign seg_2_22_lutff_0_out_9801 = net_9801;
  assign seg_2_22_lutff_5_out_9806 = net_9806;
  assign seg_2_22_neigh_op_tnl_2_4768 = seg_1_23_lutff_2_out_4768;
  assign seg_2_23_lutff_4_out_9952 = net_9952;
  assign seg_2_25_sp4_h_l_39_5472 = seg_0_25_sp4_h_r_26_5472;
  assign seg_2_26_sp4_h_l_41_5683 = seg_0_26_sp4_h_r_28_5683;
  assign seg_2_2_lutff_0_out_6825 = net_6825;
  assign seg_2_2_lutff_1_out_6826 = net_6826;
  assign seg_2_2_lutff_2_out_6827 = net_6827;
  assign seg_2_2_lutff_3_out_6828 = net_6828;
  assign seg_2_2_lutff_4_out_6829 = net_6829;
  assign seg_2_2_lutff_5_out_6830 = net_6830;
  assign seg_2_2_lutff_6_out_6831 = net_6831;
  assign seg_2_2_lutff_7_out_6832 = net_6832;
  assign seg_2_2_neigh_op_bnr_6_11235 = seg_3_1_lutff_6_out_11235;
  assign seg_2_2_neigh_op_bot_3_6676 = seg_2_1_lutff_3_out_6676;
  assign seg_2_2_neigh_op_bot_5_6678 = seg_2_1_lutff_5_out_6678;
  assign seg_2_2_neigh_op_lft_1_117 = seg_1_2_lutff_1_out_117;
  assign seg_2_2_neigh_op_lft_2_118 = seg_1_2_lutff_2_out_118;
  assign seg_2_2_neigh_op_lft_4_120 = seg_1_2_lutff_4_out_120;
  assign seg_2_2_neigh_op_lft_5_121 = seg_1_2_lutff_5_out_121;
  assign seg_2_2_neigh_op_tnl_4_455 = seg_1_3_lutff_4_out_455;
  assign seg_2_2_neigh_op_top_2_7010 = seg_2_3_lutff_2_out_7010;
  assign seg_2_2_neigh_op_top_3_7011 = seg_2_3_lutff_3_out_7011;
  assign seg_2_2_neigh_op_top_6_7014 = seg_2_3_lutff_6_out_7014;
  assign seg_2_2_sp4_h_r_0_11528 = net_11528;
  assign seg_2_2_sp4_h_r_22_7023 = net_7023;
  assign seg_2_2_sp4_h_r_41_523 = seg_1_2_sp4_h_r_28_523;
  assign seg_2_2_sp4_h_r_6_11536 = net_11536;
  assign seg_2_2_sp4_h_r_8_11538 = net_11538;
  assign seg_2_2_sp4_r_v_b_39_11543 = net_11543;
  assign seg_2_2_sp4_v_b_36_7032 = seg_1_5_sp4_r_v_b_1_7032;
  assign seg_2_2_sp4_v_b_40_7036 = net_7036;
  assign seg_2_2_sp4_v_t_36_7179 = seg_2_5_sp4_v_b_12_7179;
  assign seg_2_3_lutff_0_out_7008 = net_7008;
  assign seg_2_3_lutff_1_out_7009 = net_7009;
  assign seg_2_3_lutff_2_out_7010 = net_7010;
  assign seg_2_3_lutff_3_out_7011 = net_7011;
  assign seg_2_3_lutff_4_out_7012 = net_7012;
  assign seg_2_3_lutff_5_out_7013 = net_7013;
  assign seg_2_3_lutff_6_out_7014 = net_7014;
  assign seg_2_3_lutff_7_out_7015 = net_7015;
  assign seg_2_3_neigh_op_bot_0_6825 = seg_2_2_lutff_0_out_6825;
  assign seg_2_3_neigh_op_bot_1_6826 = seg_2_2_lutff_1_out_6826;
  assign seg_2_3_neigh_op_bot_4_6829 = seg_2_2_lutff_4_out_6829;
  assign seg_2_3_neigh_op_bot_6_6831 = seg_2_2_lutff_6_out_6831;
  assign seg_2_3_neigh_op_lft_2_453 = seg_1_3_lutff_2_out_453;
  assign seg_2_3_neigh_op_lft_4_455 = seg_1_3_lutff_4_out_455;
  assign seg_2_3_neigh_op_tnr_7_11646 = seg_3_4_lutff_7_out_11646;
  assign seg_2_3_neigh_op_top_3_7158 = seg_2_4_lutff_3_out_7158;
  assign seg_2_3_neigh_op_top_5_7160 = seg_2_4_lutff_5_out_7160;
  assign seg_2_3_sp4_h_l_38_761 = seg_1_3_sp4_h_r_38_761;
  assign seg_2_3_sp4_h_r_23_7169 = seg_1_3_sp4_h_r_10_7169;
  assign seg_2_3_sp4_r_v_b_21_11421 = net_11421;
  assign seg_2_3_sp4_r_v_b_23_11423 = net_11423;
  assign seg_2_3_sp4_v_b_5_6871 = seg_1_1_sp4_r_v_b_29_6871;
  assign seg_2_4_lutff_0_out_7155 = net_7155;
  assign seg_2_4_lutff_1_out_7156 = net_7156;
  assign seg_2_4_lutff_2_out_7157 = net_7157;
  assign seg_2_4_lutff_3_out_7158 = net_7158;
  assign seg_2_4_lutff_4_out_7159 = net_7159;
  assign seg_2_4_lutff_5_out_7160 = net_7160;
  assign seg_2_4_lutff_6_out_7161 = net_7161;
  assign seg_2_4_lutff_7_out_7162 = net_7162;
  assign seg_2_4_neigh_op_bnl_3_454 = seg_1_3_lutff_3_out_454;
  assign seg_2_4_neigh_op_bnl_5_456 = seg_1_3_lutff_5_out_456;
  assign seg_2_4_neigh_op_bnl_6_457 = seg_1_3_lutff_6_out_457;
  assign seg_2_4_neigh_op_bot_2_7010 = seg_2_3_lutff_2_out_7010;
  assign seg_2_4_neigh_op_bot_3_7011 = seg_2_3_lutff_3_out_7011;
  assign seg_2_4_neigh_op_lft_2_680 = seg_1_4_lutff_2_out_680;
  assign seg_2_4_neigh_op_lft_4_682 = seg_1_4_lutff_4_out_682;
  assign seg_2_4_neigh_op_lft_5_683 = seg_1_4_lutff_5_out_683;
  assign seg_2_4_neigh_op_lft_7_685 = seg_1_4_lutff_7_out_685;
  assign seg_2_4_neigh_op_rgt_3_11642 = seg_3_4_lutff_3_out_11642;
  assign seg_2_4_neigh_op_rgt_4_11643 = seg_3_4_lutff_4_out_11643;
  assign seg_2_4_neigh_op_rgt_6_11645 = seg_3_4_lutff_6_out_11645;
  assign seg_2_4_neigh_op_tnr_0_11762 = seg_3_5_lutff_0_out_11762;
  assign seg_2_4_neigh_op_top_6_7308 = seg_2_5_lutff_6_out_7308;
  assign seg_2_4_sp4_h_r_10_11776 = net_11776;
  assign seg_2_4_sp4_v_b_10_6891 = net_6891;
  assign seg_2_4_sp4_v_b_16_7036 = seg_2_2_sp4_v_b_40_7036;
  assign seg_2_4_sp4_v_b_8_6889 = seg_1_1_sp4_r_v_b_45_6889;
  assign seg_2_5_lutff_2_out_7304 = net_7304;
  assign seg_2_5_lutff_4_out_7306 = net_7306;
  assign seg_2_5_lutff_6_out_7308 = net_7308;
  assign seg_2_5_lutff_7_out_7309 = net_7309;
  assign seg_2_5_neigh_op_bnl_2_680 = seg_1_4_lutff_2_out_680;
  assign seg_2_5_neigh_op_lft_6_911 = seg_1_5_lutff_6_out_911;
  assign seg_2_5_neigh_op_rgt_0_11762 = seg_3_5_lutff_0_out_11762;
  assign seg_2_5_neigh_op_rgt_4_11766 = seg_3_5_lutff_4_out_11766;
  assign seg_2_5_neigh_op_rgt_6_11768 = seg_3_5_lutff_6_out_11768;
  assign seg_2_5_sp4_h_l_37_1195 = seg_0_5_sp4_h_r_24_1195;
  assign seg_2_5_sp4_h_l_41_1199 = seg_0_5_sp4_h_r_28_1199;
  assign seg_2_5_sp4_h_l_47_1206 = seg_0_5_sp4_h_r_34_1206;
  assign seg_2_5_sp4_h_r_32_1224 = net_1224;
  assign seg_2_5_sp4_h_r_5_11904 = seg_5_5_sp4_h_r_40_11904;
  assign seg_2_5_sp4_r_v_b_29_11790 = net_11790;
  assign seg_2_5_sp4_r_v_b_39_11912 = net_11912;
  assign seg_2_5_sp4_v_b_12_7179 = net_7179;
  assign seg_2_5_sp4_v_b_32_7335 = net_7335;
  assign seg_2_6_lutff_0_out_7449 = net_7449;
  assign seg_2_6_lutff_3_out_7452 = net_7452;
  assign seg_2_6_lutff_4_out_7453 = net_7453;
  assign seg_2_6_lutff_5_out_7454 = net_7454;
  assign seg_2_6_neigh_op_tnr_1_12009 = seg_3_7_lutff_1_out_12009;
  assign seg_2_6_neigh_op_tnr_4_12012 = seg_3_7_lutff_4_out_12012;
  assign seg_2_6_neigh_op_tnr_6_12014 = seg_3_7_lutff_6_out_12014;
  assign seg_2_6_neigh_op_tnr_7_12015 = seg_3_7_lutff_7_out_12015;
  assign seg_2_6_sp4_h_r_10_12022 = net_12022;
  assign seg_2_6_sp4_h_r_20_7619 = net_7619;
  assign seg_2_6_sp4_h_r_32_1430 = seg_0_6_sp4_h_r_8_1430;
  assign seg_2_6_sp4_h_r_34_1386 = net_1386;
  assign seg_2_6_sp4_r_v_b_13_11787 = net_11787;
  assign seg_2_6_sp4_r_v_b_21_11795 = net_11795;
  assign seg_2_7_lutff_0_out_7596 = net_7596;
  assign seg_2_7_lutff_3_out_7599 = net_7599;
  assign seg_2_7_lutff_4_out_7600 = net_7600;
  assign seg_2_7_lutff_6_out_7602 = net_7602;
  assign seg_2_7_lutff_7_out_7603 = net_7603;
  assign seg_2_7_neigh_op_lft_1_1337 = seg_1_7_lutff_1_out_1337;
  assign seg_2_7_sp4_h_l_45_1618 = seg_0_7_sp4_h_r_32_1618;
  assign seg_2_7_sp4_r_v_b_3_11788 = net_11788;
  assign seg_2_7_sp4_v_b_36_7767 = seg_2_9_sp4_v_b_12_7767;
  assign seg_2_7_sp4_v_b_40_7771 = seg_1_10_sp4_r_v_b_5_7771;
  assign seg_2_7_sp4_v_b_8_7335 = seg_2_5_sp4_v_b_32_7335;
  assign seg_2_7_sp4_v_t_37_7915 = seg_1_10_sp4_r_v_b_13_7915;
  assign seg_2_7_sp4_v_t_42_7920 = seg_1_11_sp4_r_v_b_7_7920;
  assign seg_2_8_lutff_2_out_7745 = net_7745;
  assign seg_2_8_lutff_5_out_7748 = net_7748;
  assign seg_2_8_lutff_6_out_7749 = net_7749;
  assign seg_2_8_lutff_7_out_7750 = net_7750;
  assign seg_2_8_neigh_op_bot_3_7599 = seg_2_7_lutff_3_out_7599;
  assign seg_2_8_neigh_op_bot_4_7600 = seg_2_7_lutff_4_out_7600;
  assign seg_2_8_neigh_op_bot_6_7602 = seg_2_7_lutff_6_out_7602;
  assign seg_2_8_neigh_op_bot_7_7603 = seg_2_7_lutff_7_out_7603;
  assign seg_2_8_neigh_op_top_6_7896 = seg_2_9_lutff_6_out_7896;
  assign seg_2_8_sp4_h_r_6_12274 = net_12274;
  assign seg_2_8_sp4_h_r_8_12276 = net_12276;
  assign seg_2_8_sp4_r_v_b_33_12163 = net_12163;
  assign seg_2_8_sp4_r_v_b_35_12165 = net_12165;
  assign seg_2_8_sp4_v_b_29_7771 = seg_1_10_sp4_r_v_b_5_7771;
  assign seg_2_8_sp4_v_b_37_7915 = seg_1_10_sp4_r_v_b_13_7915;
  assign seg_2_8_sp4_v_t_40_8065 = seg_1_10_sp4_r_v_b_29_8065;
  assign seg_2_9_lutff_0_out_7890 = net_7890;
  assign seg_2_9_lutff_1_out_7891 = net_7891;
  assign seg_2_9_lutff_2_out_7892 = net_7892;
  assign seg_2_9_lutff_4_out_7894 = net_7894;
  assign seg_2_9_lutff_5_out_7895 = net_7895;
  assign seg_2_9_lutff_6_out_7896 = net_7896;
  assign seg_2_9_neigh_op_lft_5_1758 = seg_1_9_lutff_5_out_1758;
  assign seg_2_9_neigh_op_lft_7_1760 = seg_1_9_lutff_7_out_1760;
  assign seg_2_9_neigh_op_tnl_1_1966 = seg_1_10_lutff_1_out_1966;
  assign seg_2_9_sp12_h_r_12_2012 = seg_6_9_sp12_h_r_20_2012;
  assign seg_2_9_sp4_h_r_0_12389 = seg_4_9_sp4_h_r_24_12389;
  assign seg_2_9_sp4_h_r_12_8050 = net_8050;
  assign seg_2_9_sp4_h_r_22_8052 = net_8052;
  assign seg_2_9_sp4_h_r_8_12399 = seg_4_9_sp4_h_r_32_12399;
  assign seg_2_9_sp4_r_v_b_13_12156 = net_12156;
  assign seg_2_9_sp4_r_v_b_23_12166 = net_12166;
  assign seg_2_9_sp4_r_v_b_31_12284 = net_12284;
  assign seg_2_9_sp4_r_v_b_39_12404 = net_12404;
  assign seg_2_9_sp4_v_b_12_7767 = net_7767;
  assign seg_2_9_sp4_v_b_32_7923 = seg_2_11_sp4_v_b_8_7923;
  assign seg_2_9_sp4_v_b_46_8071 = net_8071;
  assign seg_2_9_sp4_v_t_47_8219 = seg_2_13_sp4_v_b_10_8219;
  assign seg_3_10_lutff_0_out_12377 = net_12377;
  assign seg_3_10_lutff_1_out_12378 = net_12378;
  assign seg_3_10_lutff_3_out_12380 = net_12380;
  assign seg_3_10_lutff_4_out_12381 = net_12381;
  assign seg_3_10_lutff_5_out_12382 = net_12382;
  assign seg_3_10_lutff_7_out_12384 = net_12384;
  assign seg_3_10_neigh_op_top_4_12504 = seg_3_11_lutff_4_out_12504;
  assign seg_3_10_sp4_h_l_42_2248 = seg_2_10_sp4_h_r_42_2248;
  assign seg_3_10_sp4_h_r_11_16346 = seg_4_10_sp4_h_r_22_16346;
  assign seg_3_10_sp4_h_r_4_16349 = net_16349;
  assign seg_3_10_sp4_h_r_9_16354 = seg_4_10_sp4_h_r_20_16354;
  assign seg_3_10_sp4_r_v_b_29_16236 = net_16236;
  assign seg_3_10_sp4_v_b_0_12156 = seg_2_9_sp4_r_v_b_13_12156;
  assign seg_3_10_sp4_v_b_10_12166 = seg_2_9_sp4_r_v_b_23_12166;
  assign seg_3_10_sp4_v_b_11_12165 = seg_2_8_sp4_r_v_b_35_12165;
  assign seg_3_10_sp4_v_b_4_12160 = net_12160;
  assign seg_3_10_sp4_v_b_8_12164 = seg_3_8_sp4_v_b_32_12164;
  assign seg_3_10_sp4_v_b_9_12163 = seg_2_8_sp4_r_v_b_33_12163;
  assign seg_3_10_sp4_v_t_43_12654 = seg_3_14_sp4_v_b_6_12654;
  assign seg_3_11_lutff_2_out_12502 = net_12502;
  assign seg_3_11_lutff_4_out_12504 = net_12504;
  assign seg_3_11_lutff_7_out_12507 = net_12507;
  assign seg_3_11_neigh_op_lft_5_8189 = seg_2_11_lutff_5_out_8189;
  assign seg_3_11_sp4_h_l_36_2448 = seg_0_11_sp4_h_r_12_2448;
  assign seg_3_11_sp4_h_r_11_16469 = seg_6_11_sp4_h_r_46_16469;
  assign seg_3_11_sp4_h_r_3_16471 = seg_6_11_sp4_h_r_38_16471;
  assign seg_3_11_sp4_h_r_42_2489 = net_2489;
  assign seg_3_11_sp4_h_r_44_2491 = net_2491;
  assign seg_3_11_sp4_h_r_8_16476 = seg_5_11_sp4_h_r_32_16476;
  assign seg_3_11_sp4_r_v_b_1_16109 = net_16109;
  assign seg_3_11_sp4_r_v_b_27_16357 = net_16357;
  assign seg_3_11_sp4_r_v_b_29_16359 = net_16359;
  assign seg_3_11_sp4_r_v_b_33_16363 = net_16363;
  assign seg_3_11_sp4_r_v_b_3_16111 = net_16111;
  assign seg_3_11_sp4_r_v_b_7_16115 = net_16115;
  assign seg_3_11_sp4_v_b_11_12288 = seg_3_8_sp4_v_b_46_12288;
  assign seg_3_11_sp4_v_b_18_12407 = net_12407;
  assign seg_3_11_sp4_v_b_22_12411 = net_12411;
  assign seg_3_11_sp4_v_b_7_12284 = seg_2_9_sp4_r_v_b_31_12284;
  assign seg_3_12_lutff_1_out_12624 = net_12624;
  assign seg_3_12_lutff_2_out_12625 = net_12625;
  assign seg_3_12_lutff_3_out_12626 = net_12626;
  assign seg_3_12_lutff_4_out_12627 = net_12627;
  assign seg_3_12_lutff_5_out_12628 = net_12628;
  assign seg_3_12_lutff_6_out_12629 = net_12629;
  assign seg_3_12_lutff_7_out_12630 = net_12630;
  assign seg_3_12_neigh_op_bot_7_12507 = seg_3_11_lutff_7_out_12507;
  assign seg_3_12_neigh_op_rgt_2_16456 = seg_4_12_lutff_2_out_16456;
  assign seg_3_12_neigh_op_tnl_4_8482 = seg_2_13_lutff_4_out_8482;
  assign seg_3_12_neigh_op_tnl_6_8484 = seg_2_13_lutff_6_out_8484;
  assign seg_3_12_sp4_h_l_37_2657 = seg_1_12_sp4_h_r_24_2657;
  assign seg_3_12_sp4_h_l_40_2660 = seg_0_12_sp4_h_r_16_2660;
  assign seg_3_12_sp4_h_l_44_2665 = seg_0_12_sp4_h_r_20_2665;
  assign seg_3_12_sp4_h_r_10_16591 = seg_5_12_sp4_h_r_34_16591;
  assign seg_3_12_sp4_h_r_13_12758 = seg_4_12_sp4_h_r_24_12758;
  assign seg_3_12_sp4_h_r_4_16595 = seg_5_12_sp4_h_r_28_16595;
  assign seg_3_12_sp4_r_v_b_39_16604 = seg_3_14_sp4_r_v_b_15_16604;
  assign seg_3_12_sp4_v_b_11_12411 = seg_3_11_sp4_v_b_22_12411;
  assign seg_3_12_sp4_v_b_13_12525 = seg_2_10_sp4_r_v_b_37_12525;
  assign seg_3_12_sp4_v_b_2_12404 = seg_2_9_sp4_r_v_b_39_12404;
  assign seg_3_12_sp4_v_b_36_12770 = seg_3_14_sp4_v_b_12_12770;
  assign seg_3_12_sp4_v_b_7_12407 = seg_3_11_sp4_v_b_18_12407;
  assign seg_3_12_sp4_v_t_37_12894 = seg_3_14_sp4_v_b_24_12894;
  assign seg_3_12_sp4_v_t_42_12899 = seg_2_14_sp4_r_v_b_31_12899;
  assign seg_3_12_sp4_v_t_43_12900 = seg_3_16_sp4_v_b_6_12900;
  assign seg_3_12_sp4_v_t_46_12903 = seg_2_14_sp4_r_v_b_35_12903;
  assign seg_3_13_lutff_7_out_12753 = net_12753;
  assign seg_3_13_neigh_op_bnl_0_8331 = seg_2_12_lutff_0_out_8331;
  assign seg_3_13_neigh_op_bnl_1_8332 = seg_2_12_lutff_1_out_8332;
  assign seg_3_13_neigh_op_bnl_2_8333 = seg_2_12_lutff_2_out_8333;
  assign seg_3_13_neigh_op_bnl_3_8334 = seg_2_12_lutff_3_out_8334;
  assign seg_3_13_neigh_op_bnl_4_8335 = seg_2_12_lutff_4_out_8335;
  assign seg_3_13_neigh_op_bnl_5_8336 = seg_2_12_lutff_5_out_8336;
  assign seg_3_13_neigh_op_bnl_6_8337 = seg_2_12_lutff_6_out_8337;
  assign seg_3_13_neigh_op_top_5_12874 = seg_3_14_lutff_5_out_12874;
  assign seg_3_13_sp4_h_l_39_2868 = seg_1_13_sp4_h_r_26_2868;
  assign seg_3_13_sp4_h_l_41_2870 = seg_1_13_sp4_h_r_28_2870;
  assign seg_3_13_sp4_h_l_43_2872 = seg_1_13_sp4_h_r_30_2872;
  assign seg_3_13_sp4_h_r_10_16714 = net_16714;
  assign seg_3_13_sp4_h_r_12_12882 = net_12882;
  assign seg_3_13_sp4_h_r_20_12892 = net_12892;
  assign seg_3_13_sp4_h_r_22_12884 = net_12884;
  assign seg_3_13_sp4_h_r_2_16716 = net_16716;
  assign seg_3_13_sp4_h_r_8_16722 = net_16722;
  assign seg_3_13_sp4_r_v_b_31_16607 = seg_3_15_sp4_r_v_b_7_16607;
  assign seg_3_13_sp4_r_v_b_37_16725 = seg_3_15_sp4_r_v_b_13_16725;
  assign seg_3_13_sp4_r_v_b_43_16731 = seg_3_15_sp4_r_v_b_19_16731;
  assign seg_3_13_sp4_v_b_28_12775 = seg_3_15_sp4_v_b_4_12775;
  assign seg_3_13_sp4_v_b_32_12779 = seg_3_15_sp4_v_b_8_12779;
  assign seg_3_13_sp4_v_b_34_12781 = seg_3_15_sp4_v_b_10_12781;
  assign seg_3_13_sp4_v_b_38_12895 = seg_3_15_sp4_v_b_14_12895;
  assign seg_3_13_sp4_v_b_7_12530 = seg_2_11_sp4_r_v_b_31_12530;
  assign seg_3_13_sp4_v_t_36_13016 = seg_3_16_sp4_v_b_12_13016;
  assign seg_3_13_sp4_v_t_37_13017 = seg_3_17_sp4_v_b_0_13017;
  assign seg_3_14_lutff_0_out_12869 = net_12869;
  assign seg_3_14_lutff_1_out_12870 = net_12870;
  assign seg_3_14_lutff_2_out_12871 = net_12871;
  assign seg_3_14_lutff_5_out_12874 = net_12874;
  assign seg_3_14_neigh_op_bnl_0_8478 = seg_2_13_lutff_0_out_8478;
  assign seg_3_14_neigh_op_rgt_0_16700 = seg_4_14_lutff_0_out_16700;
  assign seg_3_14_neigh_op_rgt_3_16703 = seg_4_14_lutff_3_out_16703;
  assign seg_3_14_neigh_op_tnr_5_16828 = seg_4_15_lutff_5_out_16828;
  assign seg_3_14_neigh_op_top_7_12999 = seg_3_15_lutff_7_out_12999;
  assign seg_3_14_sp4_h_l_36_3092 = seg_2_14_sp4_h_r_36_3092;
  assign seg_3_14_sp4_r_v_b_15_16604 = net_16604;
  assign seg_3_14_sp4_v_b_12_12770 = net_12770;
  assign seg_3_14_sp4_v_b_24_12894 = net_12894;
  assign seg_3_14_sp4_v_b_28_12898 = seg_3_16_sp4_v_b_4_12898;
  assign seg_3_14_sp4_v_b_6_12654 = net_12654;
  assign seg_3_14_sp4_v_b_7_12653 = seg_2_12_sp4_r_v_b_31_12653;
  assign seg_3_14_sp4_v_t_45_13148 = seg_3_18_sp4_v_b_8_13148;
  assign seg_3_15_lutff_7_out_12999 = net_12999;
  assign seg_3_15_neigh_op_bnr_3_16703 = seg_4_14_lutff_3_out_16703;
  assign seg_3_15_neigh_op_lft_6_8778 = seg_2_15_lutff_6_out_8778;
  assign seg_3_15_neigh_op_rgt_2_16825 = seg_4_15_lutff_2_out_16825;
  assign seg_3_15_neigh_op_rgt_3_16826 = seg_4_15_lutff_3_out_16826;
  assign seg_3_15_neigh_op_rgt_4_16827 = seg_4_15_lutff_4_out_16827;
  assign seg_3_15_neigh_op_tnl_4_8923 = seg_2_16_lutff_4_out_8923;
  assign seg_3_15_neigh_op_tnl_5_8924 = seg_2_16_lutff_5_out_8924;
  assign seg_3_15_neigh_op_tnr_6_16952 = seg_4_16_lutff_6_out_16952;
  assign seg_3_15_neigh_op_top_0_13115 = seg_3_16_lutff_0_out_13115;
  assign seg_3_15_neigh_op_top_1_13116 = seg_3_16_lutff_1_out_13116;
  assign seg_3_15_neigh_op_top_2_13117 = seg_3_16_lutff_2_out_13117;
  assign seg_3_15_neigh_op_top_4_13119 = seg_3_16_lutff_4_out_13119;
  assign seg_3_15_neigh_op_top_5_13120 = seg_3_16_lutff_5_out_13120;
  assign seg_3_15_sp4_h_l_38_3304 = seg_0_15_sp4_h_r_14_3304;
  assign seg_3_15_sp4_h_l_40_3306 = seg_0_15_sp4_h_r_16_3306;
  assign seg_3_15_sp4_h_l_42_3308 = seg_0_15_sp4_h_r_18_3308;
  assign seg_3_15_sp4_r_v_b_13_16725 = net_16725;
  assign seg_3_15_sp4_r_v_b_19_16731 = net_16731;
  assign seg_3_15_sp4_r_v_b_7_16607 = net_16607;
  assign seg_3_15_sp4_v_b_10_12781 = net_12781;
  assign seg_3_15_sp4_v_b_14_12895 = net_12895;
  assign seg_3_15_sp4_v_b_38_13141 = seg_3_17_sp4_v_b_14_13141;
  assign seg_3_15_sp4_v_b_4_12775 = net_12775;
  assign seg_3_15_sp4_v_b_8_12779 = net_12779;
  assign seg_3_15_sp4_v_t_38_13264 = seg_3_18_sp4_v_b_14_13264;
  assign seg_3_16_lutff_0_out_13115 = net_13115;
  assign seg_3_16_lutff_1_out_13116 = net_13116;
  assign seg_3_16_lutff_2_out_13117 = net_13117;
  assign seg_3_16_lutff_4_out_13119 = net_13119;
  assign seg_3_16_lutff_5_out_13120 = net_13120;
  assign seg_3_16_lutff_7_out_13122 = net_13122;
  assign seg_3_16_neigh_op_lft_3_8922 = seg_2_16_lutff_3_out_8922;
  assign seg_3_16_neigh_op_rgt_1_16947 = seg_4_16_lutff_1_out_16947;
  assign seg_3_16_neigh_op_tnl_5_9071 = seg_2_17_lutff_5_out_9071;
  assign seg_3_16_neigh_op_top_2_13240 = seg_3_17_lutff_2_out_13240;
  assign seg_3_16_neigh_op_top_3_13241 = seg_3_17_lutff_3_out_13241;
  assign seg_3_16_neigh_op_top_4_13242 = seg_3_17_lutff_4_out_13242;
  assign seg_3_16_neigh_op_top_5_13243 = seg_3_17_lutff_5_out_13243;
  assign seg_3_16_neigh_op_top_6_13244 = seg_3_17_lutff_6_out_13244;
  assign seg_3_16_sp4_h_l_42_3514 = seg_0_16_sp4_h_r_18_3514;
  assign seg_3_16_sp4_v_b_12_13016 = net_13016;
  assign seg_3_16_sp4_v_b_4_12898 = net_12898;
  assign seg_3_16_sp4_v_b_6_12900 = net_12900;
  assign seg_3_16_sp4_v_t_39_13388 = seg_3_20_sp4_v_b_2_13388;
  assign seg_3_17_lutff_2_out_13240 = net_13240;
  assign seg_3_17_lutff_3_out_13241 = net_13241;
  assign seg_3_17_lutff_4_out_13242 = net_13242;
  assign seg_3_17_lutff_5_out_13243 = net_13243;
  assign seg_3_17_lutff_6_out_13244 = net_13244;
  assign seg_3_17_neigh_op_tnl_0_9213 = seg_2_18_lutff_0_out_9213;
  assign seg_3_17_neigh_op_tnl_1_9214 = seg_2_18_lutff_1_out_9214;
  assign seg_3_17_neigh_op_tnl_6_9219 = seg_2_18_lutff_6_out_9219;
  assign seg_3_17_neigh_op_tnl_7_9220 = seg_2_18_lutff_7_out_9220;
  assign seg_3_17_sp4_h_r_10_17206 = seg_5_17_sp4_h_r_34_17206;
  assign seg_3_17_sp4_r_v_b_29_17097 = seg_3_19_sp4_r_v_b_5_17097;
  assign seg_3_17_sp4_v_b_0_13017 = net_13017;
  assign seg_3_17_sp4_v_b_14_13141 = net_13141;
  assign seg_3_17_sp4_v_t_47_13519 = seg_3_21_sp4_v_b_10_13519;
  assign seg_3_18_neigh_op_tnl_4_9364 = seg_2_19_lutff_4_out_9364;
  assign seg_3_18_neigh_op_top_5_13489 = seg_3_19_lutff_5_out_13489;
  assign seg_3_18_sp4_r_v_b_11_16980 = net_16980;
  assign seg_3_18_sp4_r_v_b_13_17094 = net_17094;
  assign seg_3_18_sp4_r_v_b_1_16970 = net_16970;
  assign seg_3_18_sp4_v_b_14_13264 = net_13264;
  assign seg_3_18_sp4_v_b_8_13148 = net_13148;
  assign seg_3_18_sp4_v_t_36_13631 = seg_3_21_sp4_v_b_12_13631;
  assign seg_3_19_lutff_5_out_13489 = net_13489;
  assign seg_3_19_neigh_op_lft_0_9360 = seg_2_19_lutff_0_out_9360;
  assign seg_3_19_neigh_op_tnl_1_9508 = seg_2_20_lutff_1_out_9508;
  assign seg_3_19_sp4_r_v_b_5_17097 = net_17097;
  assign seg_3_1_lutff_0_out_11229 = net_11229;
  assign seg_3_1_lutff_1_out_11230 = net_11230;
  assign seg_3_1_lutff_2_out_11231 = net_11231;
  assign seg_3_1_lutff_3_out_11232 = net_11232;
  assign seg_3_1_lutff_6_out_11235 = net_11235;
  assign seg_3_1_lutff_7_out_11236 = net_11236;
  assign seg_3_1_neigh_op_rgt_0_15060 = seg_4_1_lutff_0_out_15060;
  assign seg_3_1_neigh_op_rgt_3_15063 = seg_4_1_lutff_3_out_15063;
  assign seg_3_1_neigh_op_rgt_5_15065 = seg_4_1_lutff_5_out_15065;
  assign seg_3_1_neigh_op_rgt_6_15066 = seg_4_1_lutff_6_out_15066;
  assign seg_3_1_neigh_op_rgt_7_15067 = seg_4_1_lutff_7_out_15067;
  assign seg_3_1_neigh_op_tnl_3_6828 = seg_2_2_lutff_3_out_6828;
  assign seg_3_1_neigh_op_tnr_6_15194 = seg_4_2_lutff_6_out_15194;
  assign seg_3_1_sp4_h_r_12_11370 = net_11370;
  assign seg_3_1_sp4_h_r_14_11374 = net_11374;
  assign seg_3_1_sp4_h_r_18_11378 = net_11378;
  assign seg_3_1_sp4_h_r_20_11380 = net_11380;
  assign seg_3_1_sp4_h_r_44_250 = net_250;
  assign seg_3_1_sp4_h_r_6_15208 = net_15208;
  assign seg_3_1_sp4_r_v_b_29_15234 = net_15234;
  assign seg_3_1_sp4_v_b_41_11417 = seg_3_4_sp4_v_b_4_11417;
  assign seg_3_1_sp4_v_t_37_11541 = seg_3_5_sp4_v_b_0_11541;
  assign seg_3_1_sp4_v_t_44_11548 = seg_3_4_sp4_v_b_20_11548;
  assign seg_3_20_sp4_v_b_2_13388 = net_13388;
  assign seg_3_21_neigh_op_top_3_13856 = seg_3_22_lutff_3_out_13856;
  assign seg_3_21_sp4_v_b_10_13519 = net_13519;
  assign seg_3_21_sp4_v_b_12_13631 = net_13631;
  assign seg_3_22_lutff_3_out_13856 = net_13856;
  assign seg_3_22_neigh_op_tnl_4_9952 = seg_2_23_lutff_4_out_9952;
  assign seg_3_24_sp4_h_l_46_5260 = seg_0_24_sp4_h_r_22_5260;
  assign seg_3_2_lutff_0_out_11357 = net_11357;
  assign seg_3_2_lutff_1_out_11358 = net_11358;
  assign seg_3_2_lutff_2_out_11359 = net_11359;
  assign seg_3_2_lutff_3_out_11360 = net_11360;
  assign seg_3_2_lutff_4_out_11361 = net_11361;
  assign seg_3_2_lutff_5_out_11362 = net_11362;
  assign seg_3_2_lutff_6_out_11363 = net_11363;
  assign seg_3_2_lutff_7_out_11364 = net_11364;
  assign seg_3_2_neigh_op_bnr_3_15063 = seg_4_1_lutff_3_out_15063;
  assign seg_3_2_neigh_op_rgt_1_15189 = seg_4_2_lutff_1_out_15189;
  assign seg_3_2_neigh_op_rgt_4_15192 = seg_4_2_lutff_4_out_15192;
  assign seg_3_2_neigh_op_rgt_5_15193 = seg_4_2_lutff_5_out_15193;
  assign seg_3_2_neigh_op_top_0_11516 = seg_3_3_lutff_0_out_11516;
  assign seg_3_2_sp4_h_r_4_15365 = net_15365;
  assign seg_3_2_sp4_h_r_8_15369 = net_15369;
  assign seg_3_2_sp4_r_v_b_13_15229 = net_15229;
  assign seg_3_2_sp4_r_v_b_24_15243 = seg_4_4_sp4_v_b_0_15243;
  assign seg_3_2_sp4_r_v_b_29_15247 = seg_3_4_sp4_r_v_b_5_15247;
  assign seg_3_2_sp4_r_v_b_31_15249 = net_15249;
  assign seg_3_2_sp4_v_t_41_11668 = seg_3_4_sp4_v_b_28_11668;
  assign seg_3_3_lutff_0_out_11516 = net_11516;
  assign seg_3_3_lutff_1_out_11517 = net_11517;
  assign seg_3_3_lutff_2_out_11518 = net_11518;
  assign seg_3_3_lutff_3_out_11519 = net_11519;
  assign seg_3_3_lutff_4_out_11520 = net_11520;
  assign seg_3_3_lutff_5_out_11521 = net_11521;
  assign seg_3_3_lutff_6_out_11522 = net_11522;
  assign seg_3_3_lutff_7_out_11523 = net_11523;
  assign seg_3_3_neigh_op_bot_6_11363 = seg_3_2_lutff_6_out_11363;
  assign seg_3_3_neigh_op_rgt_0_15347 = seg_4_3_lutff_0_out_15347;
  assign seg_3_3_neigh_op_rgt_2_15349 = seg_4_3_lutff_2_out_15349;
  assign seg_3_3_neigh_op_rgt_3_15350 = seg_4_3_lutff_3_out_15350;
  assign seg_3_3_neigh_op_rgt_4_15351 = seg_4_3_lutff_4_out_15351;
  assign seg_3_3_neigh_op_tnr_0_15470 = seg_4_4_lutff_0_out_15470;
  assign seg_3_3_neigh_op_tnr_3_15473 = seg_4_4_lutff_3_out_15473;
  assign seg_3_3_neigh_op_top_2_11641 = seg_3_4_lutff_2_out_11641;
  assign seg_3_3_sp4_h_r_4_15488 = net_15488;
  assign seg_3_3_sp4_h_r_6_15490 = net_15490;
  assign seg_3_3_sp4_r_v_b_14_15244 = seg_4_1_sp4_v_b_38_15244;
  assign seg_3_3_sp4_v_b_40_11667 = net_11667;
  assign seg_3_3_sp4_v_t_40_11790 = seg_2_5_sp4_r_v_b_29_11790;
  assign seg_3_4_lutff_0_out_11639 = net_11639;
  assign seg_3_4_lutff_2_out_11641 = net_11641;
  assign seg_3_4_lutff_3_out_11642 = net_11642;
  assign seg_3_4_lutff_4_out_11643 = net_11643;
  assign seg_3_4_lutff_5_out_11644 = net_11644;
  assign seg_3_4_lutff_6_out_11645 = net_11645;
  assign seg_3_4_lutff_7_out_11646 = net_11646;
  assign seg_3_4_neigh_op_bnl_1_7009 = seg_2_3_lutff_1_out_7009;
  assign seg_3_4_neigh_op_lft_5_7160 = seg_2_4_lutff_5_out_7160;
  assign seg_3_4_neigh_op_lft_6_7161 = seg_2_4_lutff_6_out_7161;
  assign seg_3_4_neigh_op_lft_7_7162 = seg_2_4_lutff_7_out_7162;
  assign seg_3_4_neigh_op_rgt_0_15470 = seg_4_4_lutff_0_out_15470;
  assign seg_3_4_neigh_op_rgt_3_15473 = seg_4_4_lutff_3_out_15473;
  assign seg_3_4_neigh_op_top_0_11762 = seg_3_5_lutff_0_out_11762;
  assign seg_3_4_sp4_h_r_11_15608 = seg_6_4_sp4_h_r_46_15608;
  assign seg_3_4_sp4_h_r_12_11775 = net_11775;
  assign seg_3_4_sp4_h_r_1_15606 = seg_6_4_sp4_h_r_36_15606;
  assign seg_3_4_sp4_r_v_b_1_15242 = net_15242;
  assign seg_3_4_sp4_r_v_b_5_15247 = net_15247;
  assign seg_3_4_sp4_v_b_10_11423 = seg_2_3_sp4_r_v_b_23_11423;
  assign seg_3_4_sp4_v_b_15_11543 = seg_2_2_sp4_r_v_b_39_11543;
  assign seg_3_4_sp4_v_b_20_11548 = net_11548;
  assign seg_3_4_sp4_v_b_28_11668 = net_11668;
  assign seg_3_4_sp4_v_b_32_11672 = net_11672;
  assign seg_3_4_sp4_v_b_4_11417 = net_11417;
  assign seg_3_4_sp4_v_b_8_11421 = seg_2_3_sp4_r_v_b_21_11421;
  assign seg_3_4_sp4_v_t_39_11912 = seg_2_5_sp4_r_v_b_39_11912;
  assign seg_3_5_lutff_0_out_11762 = net_11762;
  assign seg_3_5_lutff_2_out_11764 = net_11764;
  assign seg_3_5_lutff_4_out_11766 = net_11766;
  assign seg_3_5_lutff_6_out_11768 = net_11768;
  assign seg_3_5_neigh_op_bot_0_11639 = seg_3_4_lutff_0_out_11639;
  assign seg_3_5_neigh_op_rgt_3_15596 = seg_4_5_lutff_3_out_15596;
  assign seg_3_5_neigh_op_tnl_5_7454 = seg_2_6_lutff_5_out_7454;
  assign seg_3_5_sp4_h_l_38_1184 = seg_0_5_sp4_h_r_14_1184;
  assign seg_3_5_sp4_h_r_10_15730 = seg_5_5_sp4_h_r_34_15730;
  assign seg_3_5_sp4_h_r_12_11898 = seg_5_5_sp4_h_r_36_11898;
  assign seg_3_5_sp4_h_r_14_11902 = seg_5_5_sp4_h_r_38_11902;
  assign seg_3_5_sp4_h_r_26_7465 = net_7465;
  assign seg_3_5_sp4_h_r_30_7469 = net_7469;
  assign seg_3_5_sp4_h_r_32_7471 = net_7471;
  assign seg_3_5_sp4_h_r_34_7463 = net_7463;
  assign seg_3_5_sp4_r_v_b_33_15625 = net_15625;
  assign seg_3_5_sp4_v_b_0_11541 = net_11541;
  assign seg_3_6_lutff_0_out_11885 = net_11885;
  assign seg_3_6_lutff_1_out_11886 = net_11886;
  assign seg_3_6_lutff_5_out_11890 = net_11890;
  assign seg_3_6_lutff_7_out_11892 = net_11892;
  assign seg_3_6_neigh_op_bnr_5_15598 = seg_4_5_lutff_5_out_15598;
  assign seg_3_6_neigh_op_rgt_0_15716 = seg_4_6_lutff_0_out_15716;
  assign seg_3_6_sp4_h_r_12_12021 = net_12021;
  assign seg_3_6_sp4_h_r_8_15861 = net_15861;
  assign seg_3_6_sp4_v_b_22_11796 = net_11796;
  assign seg_3_6_sp4_v_b_5_11667 = seg_3_3_sp4_v_b_40_11667;
  assign seg_3_6_sp4_v_b_8_11672 = seg_3_4_sp4_v_b_32_11672;
  assign seg_3_6_sp4_v_t_41_12160 = seg_3_10_sp4_v_b_4_12160;
  assign seg_3_6_sp4_v_t_47_12166 = seg_2_9_sp4_r_v_b_23_12166;
  assign seg_3_7_lutff_1_out_12009 = net_12009;
  assign seg_3_7_lutff_4_out_12012 = net_12012;
  assign seg_3_7_lutff_6_out_12014 = net_12014;
  assign seg_3_7_lutff_7_out_12015 = net_12015;
  assign seg_3_7_neigh_op_bnr_1_15717 = seg_4_6_lutff_1_out_15717;
  assign seg_3_7_neigh_op_bnr_2_15718 = seg_4_6_lutff_2_out_15718;
  assign seg_3_7_neigh_op_bnr_3_15719 = seg_4_6_lutff_3_out_15719;
  assign seg_3_7_neigh_op_bnr_5_15721 = seg_4_6_lutff_5_out_15721;
  assign seg_3_7_neigh_op_bnr_6_15722 = seg_4_6_lutff_6_out_15722;
  assign seg_3_7_sp4_h_l_38_1598 = seg_0_7_sp4_h_r_14_1598;
  assign seg_3_7_sp4_h_r_26_7759 = net_7759;
  assign seg_3_7_sp4_v_b_0_11787 = seg_2_6_sp4_r_v_b_13_11787;
  assign seg_3_7_sp4_v_b_11_11796 = seg_3_6_sp4_v_b_22_11796;
  assign seg_3_7_sp4_v_b_20_11917 = net_11917;
  assign seg_3_7_sp4_v_b_22_11919 = net_11919;
  assign seg_3_7_sp4_v_b_3_11788 = seg_2_7_sp4_r_v_b_3_11788;
  assign seg_3_7_sp4_v_b_8_11795 = seg_2_6_sp4_r_v_b_21_11795;
  assign seg_3_8_lutff_4_out_12135 = net_12135;
  assign seg_3_8_neigh_op_tnl_1_7891 = seg_2_9_lutff_1_out_7891;
  assign seg_3_8_neigh_op_tnl_4_7894 = seg_2_9_lutff_4_out_7894;
  assign seg_3_8_sp4_h_l_36_1805 = seg_0_8_sp4_h_r_12_1805;
  assign seg_3_8_sp4_h_l_44_1814 = seg_0_8_sp4_h_r_20_1814;
  assign seg_3_8_sp4_h_r_20_12277 = net_12277;
  assign seg_3_8_sp4_v_b_11_11919 = seg_3_7_sp4_v_b_22_11919;
  assign seg_3_8_sp4_v_b_32_12164 = net_12164;
  assign seg_3_8_sp4_v_b_46_12288 = net_12288;
  assign seg_3_8_sp4_v_b_9_11917 = seg_3_7_sp4_v_b_20_11917;
  assign seg_3_9_lutff_1_out_12255 = net_12255;
  assign seg_3_9_lutff_2_out_12256 = net_12256;
  assign seg_3_9_lutff_3_out_12257 = net_12257;
  assign seg_3_9_lutff_4_out_12258 = net_12258;
  assign seg_3_9_lutff_5_out_12259 = net_12259;
  assign seg_3_9_lutff_6_out_12260 = net_12260;
  assign seg_3_9_lutff_7_out_12261 = net_12261;
  assign seg_3_9_neigh_op_lft_1_7891 = seg_2_9_lutff_1_out_7891;
  assign seg_3_9_neigh_op_lft_4_7894 = seg_2_9_lutff_4_out_7894;
  assign seg_3_9_neigh_op_lft_5_7895 = seg_2_9_lutff_5_out_7895;
  assign seg_3_9_neigh_op_tnl_0_8037 = seg_2_10_lutff_0_out_8037;
  assign seg_3_9_neigh_op_tnl_6_8043 = seg_2_10_lutff_6_out_8043;
  assign seg_3_9_neigh_op_tnl_7_8044 = seg_2_10_lutff_7_out_8044;
  assign seg_3_9_neigh_op_top_0_12377 = seg_3_10_lutff_0_out_12377;
  assign seg_3_9_neigh_op_top_1_12378 = seg_3_10_lutff_1_out_12378;
  assign seg_3_9_neigh_op_top_3_12380 = seg_3_10_lutff_3_out_12380;
  assign seg_3_9_neigh_op_top_4_12381 = seg_3_10_lutff_4_out_12381;
  assign seg_3_9_neigh_op_top_7_12384 = seg_3_10_lutff_7_out_12384;
  assign seg_3_9_sp4_h_r_11_16223 = seg_4_9_sp4_h_r_22_16223;
  assign seg_3_9_sp4_h_r_3_16225 = seg_4_9_sp4_h_r_14_16225;
  assign seg_3_9_sp4_h_r_5_16227 = seg_6_9_sp4_h_r_40_16227;
  assign seg_3_9_sp4_h_r_9_16231 = seg_4_9_sp4_h_r_20_16231;
  assign seg_3_9_sp4_v_t_46_12534 = seg_2_13_sp4_r_v_b_11_12534;
  assign seg_4_0_span4_horz_r_0_18923 = seg_6_0_span4_horz_r_8_18923;
  assign seg_4_10_neigh_op_bnl_7_12261 = seg_3_9_lutff_7_out_12261;
  assign seg_4_10_sp4_h_l_36_2239 = seg_1_10_sp4_h_r_12_2239;
  assign seg_4_10_sp4_h_r_20_16354 = net_16354;
  assign seg_4_10_sp4_h_r_22_16346 = net_16346;
  assign seg_4_10_sp4_h_r_26_12516 = net_12516;
  assign seg_4_10_sp4_h_r_5_20181 = seg_5_10_sp4_h_r_16_20181;
  assign seg_4_10_sp4_r_v_b_47_20197 = net_20197;
  assign seg_4_10_sp4_v_b_24_16233 = net_16233;
  assign seg_4_10_sp4_v_b_28_16237 = net_16237;
  assign seg_4_10_sp4_v_b_32_16241 = net_16241;
  assign seg_4_10_sp4_v_b_34_16243 = net_16243;
  assign seg_4_11_sp4_h_l_37_2444 = seg_0_11_sp4_h_r_0_2444;
  assign seg_4_11_sp4_h_l_39_2456 = seg_0_11_sp4_h_r_2_2456;
  assign seg_4_11_sp4_h_l_41_2478 = seg_0_11_sp4_h_r_4_2478;
  assign seg_4_11_sp4_h_l_43_2488 = seg_0_11_sp4_h_r_6_2488;
  assign seg_4_11_sp4_h_l_45_2490 = seg_0_11_sp4_h_r_8_2490;
  assign seg_4_11_sp4_h_l_47_2446 = seg_0_11_sp4_h_r_10_2446;
  assign seg_4_11_sp4_h_r_20_16477 = seg_6_11_sp4_h_r_44_16477;
  assign seg_4_11_sp4_h_r_44_8354 = net_8354;
  assign seg_4_11_sp4_r_v_b_25_20186 = net_20186;
  assign seg_4_11_sp4_r_v_b_43_20316 = net_20316;
  assign seg_4_11_sp4_v_b_22_16242 = net_16242;
  assign seg_4_11_sp4_v_b_28_16360 = net_16360;
  assign seg_4_11_sp4_v_b_30_16362 = net_16362;
  assign seg_4_11_sp4_v_b_32_16364 = net_16364;
  assign seg_4_11_sp4_v_b_34_16366 = net_16366;
  assign seg_4_11_sp4_v_b_36_16478 = net_16478;
  assign seg_4_11_sp4_v_b_6_16116 = net_16116;
  assign seg_4_11_sp4_v_b_8_16118 = net_16118;
  assign seg_4_12_lutff_2_out_16456 = net_16456;
  assign seg_4_12_neigh_op_tnr_0_20408 = seg_5_13_lutff_0_out_20408;
  assign seg_4_12_neigh_op_tnr_2_20410 = seg_5_13_lutff_2_out_20410;
  assign seg_4_12_sp4_h_r_10_20422 = seg_6_12_sp4_h_r_34_20422;
  assign seg_4_12_sp4_h_r_18_16598 = net_16598;
  assign seg_4_12_sp4_h_r_24_12758 = net_12758;
  assign seg_4_12_sp4_h_r_4_20426 = seg_6_12_sp4_h_r_28_20426;
  assign seg_4_12_sp4_r_v_b_27_20311 = seg_4_14_sp4_r_v_b_3_20311;
  assign seg_4_12_sp4_r_v_b_39_20435 = net_20435;
  assign seg_4_12_sp4_v_b_0_16233 = seg_4_10_sp4_v_b_24_16233;
  assign seg_4_12_sp4_v_b_10_16243 = seg_4_10_sp4_v_b_34_16243;
  assign seg_4_12_sp4_v_b_11_16242 = seg_4_11_sp4_v_b_22_16242;
  assign seg_4_12_sp4_v_b_26_16481 = net_16481;
  assign seg_4_12_sp4_v_b_32_16487 = net_16487;
  assign seg_4_12_sp4_v_b_38_16603 = seg_4_14_sp4_v_b_14_16603;
  assign seg_4_12_sp4_v_b_46_16611 = net_16611;
  assign seg_4_12_sp4_v_b_4_16237 = seg_4_10_sp4_v_b_28_16237;
  assign seg_4_12_sp4_v_b_8_16241 = seg_4_10_sp4_v_b_32_16241;
  assign seg_4_13_sp4_h_l_37_2861 = seg_0_13_sp4_h_r_0_2861;
  assign seg_4_13_sp4_h_l_39_2873 = seg_2_13_sp4_h_r_26_2873;
  assign seg_4_13_sp4_h_l_46_2864 = seg_1_13_sp4_h_r_22_2864;
  assign seg_4_13_sp4_h_r_14_16717 = net_16717;
  assign seg_4_13_sp4_h_r_28_12887 = seg_2_13_sp4_h_r_4_12887;
  assign seg_4_13_sp4_h_r_30_12889 = seg_2_13_sp4_h_r_6_12889;
  assign seg_4_13_sp4_h_r_37_8637 = seg_1_13_sp4_h_r_0_8637;
  assign seg_4_13_sp4_h_r_39_8641 = seg_1_13_sp4_h_r_2_8641;
  assign seg_4_13_sp4_h_r_41_8643 = seg_1_13_sp4_h_r_4_8643;
  assign seg_4_13_sp4_h_r_45_8647 = seg_1_13_sp4_h_r_8_8647;
  assign seg_4_13_sp4_h_r_7_20552 = seg_5_13_sp4_h_r_18_20552;
  assign seg_4_13_sp4_r_v_b_19_20316 = seg_4_11_sp4_r_v_b_43_20316;
  assign seg_4_13_sp4_v_b_10_16366 = seg_4_11_sp4_v_b_34_16366;
  assign seg_4_13_sp4_v_b_12_16478 = seg_4_11_sp4_v_b_36_16478;
  assign seg_4_13_sp4_v_b_3_16357 = seg_3_11_sp4_r_v_b_27_16357;
  assign seg_4_13_sp4_v_b_4_16360 = seg_4_11_sp4_v_b_28_16360;
  assign seg_4_13_sp4_v_b_5_16359 = seg_3_11_sp4_r_v_b_29_16359;
  assign seg_4_13_sp4_v_b_6_16362 = seg_4_11_sp4_v_b_30_16362;
  assign seg_4_13_sp4_v_b_8_16364 = seg_4_11_sp4_v_b_32_16364;
  assign seg_4_13_sp4_v_b_9_16363 = seg_3_11_sp4_r_v_b_33_16363;
  assign seg_4_14_lutff_0_out_16700 = net_16700;
  assign seg_4_14_lutff_3_out_16703 = net_16703;
  assign seg_4_14_lutff_4_out_16704 = net_16704;
  assign seg_4_14_lutff_5_out_16705 = net_16705;
  assign seg_4_14_lutff_6_out_16706 = net_16706;
  assign seg_4_14_sp4_h_r_34_13006 = seg_2_14_sp4_h_r_10_13006;
  assign seg_4_14_sp4_r_v_b_3_20311 = net_20311;
  assign seg_4_14_sp4_v_b_14_16603 = net_16603;
  assign seg_4_14_sp4_v_b_2_16481 = seg_4_12_sp4_v_b_26_16481;
  assign seg_4_14_sp4_v_b_8_16487 = seg_4_12_sp4_v_b_32_16487;
  assign seg_4_14_sp4_v_t_36_16970 = seg_3_18_sp4_r_v_b_1_16970;
  assign seg_4_14_sp4_v_t_43_16977 = seg_4_18_sp4_v_b_6_16977;
  assign seg_4_14_sp4_v_t_46_16980 = seg_3_18_sp4_r_v_b_11_16980;
  assign seg_4_15_lutff_0_out_16823 = net_16823;
  assign seg_4_15_lutff_1_out_16824 = net_16824;
  assign seg_4_15_lutff_2_out_16825 = net_16825;
  assign seg_4_15_lutff_3_out_16826 = net_16826;
  assign seg_4_15_lutff_4_out_16827 = net_16827;
  assign seg_4_15_lutff_5_out_16828 = net_16828;
  assign seg_4_15_lutff_6_out_16829 = net_16829;
  assign seg_4_15_lutff_7_out_16830 = net_16830;
  assign seg_4_15_neigh_op_rgt_4_20658 = seg_5_15_lutff_4_out_20658;
  assign seg_4_15_sp4_h_l_45_3344 = seg_0_15_sp4_h_r_8_3344;
  assign seg_4_15_sp4_h_l_47_3300 = seg_0_15_sp4_h_r_10_3300;
  assign seg_4_15_sp4_h_r_34_13129 = seg_2_15_sp4_h_r_10_13129;
  assign seg_4_15_sp4_h_r_38_8936 = seg_2_15_sp4_h_r_14_8936;
  assign seg_4_15_sp4_v_b_11_16611 = seg_4_12_sp4_v_b_46_16611;
  assign seg_4_15_sp4_v_t_37_17094 = seg_3_18_sp4_r_v_b_13_17094;
  assign seg_4_16_lutff_0_out_16946 = net_16946;
  assign seg_4_16_lutff_1_out_16947 = net_16947;
  assign seg_4_16_lutff_4_out_16950 = net_16950;
  assign seg_4_16_lutff_5_out_16951 = net_16951;
  assign seg_4_16_lutff_6_out_16952 = net_16952;
  assign seg_4_16_lutff_7_out_16953 = net_16953;
  assign seg_4_16_sp4_h_r_39_9082 = seg_1_16_sp4_h_r_2_9082;
  assign seg_4_16_sp4_v_t_38_17218 = seg_4_19_sp4_v_b_14_17218;
  assign seg_4_16_sp4_v_t_40_17220 = seg_4_19_sp4_v_b_16_17220;
  assign seg_4_17_lutff_1_out_17070 = net_17070;
  assign seg_4_17_lutff_3_out_17072 = net_17072;
  assign seg_4_17_lutff_5_out_17074 = net_17074;
  assign seg_4_17_sp4_h_l_41_3746 = seg_0_17_sp4_h_r_4_3746;
  assign seg_4_17_sp4_h_l_45_3758 = seg_0_17_sp4_h_r_8_3758;
  assign seg_4_17_sp4_h_r_0_21035 = net_21035;
  assign seg_4_17_sp4_h_r_11_21038 = seg_7_17_sp4_h_r_46_21038;
  assign seg_4_17_sp4_h_r_12_17205 = net_17205;
  assign seg_4_17_sp4_h_r_8_21045 = net_21045;
  assign seg_4_17_sp4_r_v_b_31_20930 = net_20930;
  assign seg_4_18_sp4_h_l_43_3965 = seg_0_18_sp4_h_r_6_3965;
  assign seg_4_18_sp4_v_b_6_16977 = net_16977;
  assign seg_4_19_lutff_6_out_17321 = net_17321;
  assign seg_4_19_neigh_op_top_5_17443 = seg_4_20_lutff_5_out_17443;
  assign seg_4_19_sp12_v_t_23_21280 = seg_4_31_span12_vert_0_21280;
  assign seg_4_19_sp4_v_b_14_17218 = net_17218;
  assign seg_4_19_sp4_v_b_16_17220 = net_17220;
  assign seg_4_19_sp4_v_t_36_17585 = seg_4_22_sp4_v_b_12_17585;
  assign seg_4_1_lutff_0_out_15060 = net_15060;
  assign seg_4_1_lutff_2_out_15062 = net_15062;
  assign seg_4_1_lutff_3_out_15063 = net_15063;
  assign seg_4_1_lutff_4_out_15064 = net_15064;
  assign seg_4_1_lutff_5_out_15065 = net_15065;
  assign seg_4_1_lutff_6_out_15066 = net_15066;
  assign seg_4_1_lutff_7_out_15067 = net_15067;
  assign seg_4_1_neigh_op_lft_2_11231 = seg_3_1_lutff_2_out_11231;
  assign seg_4_1_neigh_op_lft_3_11232 = seg_3_1_lutff_3_out_11232;
  assign seg_4_1_neigh_op_lft_7_11236 = seg_3_1_lutff_7_out_11236;
  assign seg_4_1_neigh_op_rgt_3_18894 = seg_5_1_lutff_3_out_18894;
  assign seg_4_1_neigh_op_top_2_15190 = seg_4_2_lutff_2_out_15190;
  assign seg_4_1_neigh_op_top_3_15191 = seg_4_2_lutff_3_out_15191;
  assign seg_4_1_neigh_op_top_7_15195 = seg_4_2_lutff_7_out_15195;
  assign seg_4_1_sp4_r_v_b_39_19076 = net_19076;
  assign seg_4_1_sp4_r_v_b_41_19079 = net_19079;
  assign seg_4_1_sp4_r_v_b_43_19081 = net_19081;
  assign seg_4_1_sp4_v_b_37_15243 = seg_4_4_sp4_v_b_0_15243;
  assign seg_4_1_sp4_v_b_38_15244 = net_15244;
  assign seg_4_1_sp4_v_b_40_15247 = seg_3_4_sp4_r_v_b_5_15247;
  assign seg_4_1_sp4_v_b_43_15250 = seg_4_4_sp4_v_b_6_15250;
  assign seg_4_20_lutff_4_out_17442 = net_17442;
  assign seg_4_20_lutff_5_out_17443 = net_17443;
  assign seg_4_22_sp4_v_b_12_17585 = net_17585;
  assign seg_4_23_sp4_h_l_37_5039 = seg_0_23_sp4_h_r_0_5039;
  assign seg_4_25_sp4_h_l_37_5453 = seg_0_25_sp4_h_r_0_5453;
  assign seg_4_25_sp4_h_l_43_5497 = seg_0_25_sp4_h_r_6_5497;
  assign seg_4_25_sp4_h_l_45_5499 = seg_0_25_sp4_h_r_8_5499;
  assign seg_4_2_lutff_1_out_15189 = net_15189;
  assign seg_4_2_lutff_2_out_15190 = net_15190;
  assign seg_4_2_lutff_3_out_15191 = net_15191;
  assign seg_4_2_lutff_4_out_15192 = net_15192;
  assign seg_4_2_lutff_5_out_15193 = net_15193;
  assign seg_4_2_lutff_6_out_15194 = net_15194;
  assign seg_4_2_lutff_7_out_15195 = net_15195;
  assign seg_4_2_neigh_op_bnl_1_11230 = seg_3_1_lutff_1_out_11230;
  assign seg_4_2_neigh_op_bnl_2_11231 = seg_3_1_lutff_2_out_11231;
  assign seg_4_2_neigh_op_bnl_3_11232 = seg_3_1_lutff_3_out_11232;
  assign seg_4_2_neigh_op_bnl_7_11236 = seg_3_1_lutff_7_out_11236;
  assign seg_4_2_neigh_op_lft_2_11359 = seg_3_2_lutff_2_out_11359;
  assign seg_4_2_neigh_op_lft_4_11361 = seg_3_2_lutff_4_out_11361;
  assign seg_4_2_neigh_op_lft_7_11364 = seg_3_2_lutff_7_out_11364;
  assign seg_4_2_neigh_op_top_6_15353 = seg_4_3_lutff_6_out_15353;
  assign seg_4_2_sp4_v_b_30_15250 = seg_4_4_sp4_v_b_6_15250;
  assign seg_4_31_span12_vert_0_21280 = net_21280;
  assign seg_4_3_lutff_0_out_15347 = net_15347;
  assign seg_4_3_lutff_1_out_15348 = net_15348;
  assign seg_4_3_lutff_2_out_15349 = net_15349;
  assign seg_4_3_lutff_3_out_15350 = net_15350;
  assign seg_4_3_lutff_4_out_15351 = net_15351;
  assign seg_4_3_lutff_5_out_15352 = net_15352;
  assign seg_4_3_lutff_6_out_15353 = net_15353;
  assign seg_4_3_lutff_7_out_15354 = net_15354;
  assign seg_4_3_neigh_op_bnl_6_11363 = seg_3_2_lutff_6_out_11363;
  assign seg_4_3_neigh_op_lft_2_11518 = seg_3_3_lutff_2_out_11518;
  assign seg_4_3_neigh_op_lft_3_11519 = seg_3_3_lutff_3_out_11519;
  assign seg_4_3_neigh_op_lft_4_11520 = seg_3_3_lutff_4_out_11520;
  assign seg_4_3_neigh_op_tnl_2_11641 = seg_3_4_lutff_2_out_11641;
  assign seg_4_3_neigh_op_top_3_15473 = seg_4_4_lutff_3_out_15473;
  assign seg_4_3_neigh_op_top_6_15476 = seg_4_4_lutff_6_out_15476;
  assign seg_4_3_sp4_h_l_44_788 = seg_1_3_sp4_h_r_20_788;
  assign seg_4_3_sp4_h_r_42_7176 = net_7176;
  assign seg_4_3_sp4_r_v_b_15_19076 = seg_4_1_sp4_r_v_b_39_19076;
  assign seg_4_3_sp4_v_b_0_15229 = seg_3_2_sp4_r_v_b_13_15229;
  assign seg_4_3_sp4_v_b_5_15234 = seg_3_1_sp4_r_v_b_29_15234;
  assign seg_4_3_sp4_v_t_41_15622 = seg_4_5_sp4_v_b_28_15622;
  assign seg_4_3_sp4_v_t_44_15625 = seg_3_5_sp4_r_v_b_33_15625;
  assign seg_4_4_lutff_0_out_15470 = net_15470;
  assign seg_4_4_lutff_3_out_15473 = net_15473;
  assign seg_4_4_lutff_4_out_15474 = net_15474;
  assign seg_4_4_lutff_6_out_15476 = net_15476;
  assign seg_4_4_neigh_op_bot_6_15353 = seg_4_3_lutff_6_out_15353;
  assign seg_4_4_neigh_op_lft_2_11641 = seg_3_4_lutff_2_out_11641;
  assign seg_4_4_neigh_op_tnl_2_11764 = seg_3_5_lutff_2_out_11764;
  assign seg_4_4_sp4_h_r_26_11778 = net_11778;
  assign seg_4_4_sp4_h_r_2_19440 = net_19440;
  assign seg_4_4_sp4_h_r_4_19442 = net_19442;
  assign seg_4_4_sp4_h_r_7_19445 = seg_7_4_sp4_h_r_42_19445;
  assign seg_4_4_sp4_r_v_b_4_19079 = seg_4_1_sp4_r_v_b_41_19079;
  assign seg_4_4_sp4_r_v_b_7_19080 = net_19080;
  assign seg_4_4_sp4_v_b_0_15243 = net_15243;
  assign seg_4_4_sp4_v_b_1_15242 = seg_3_4_sp4_r_v_b_1_15242;
  assign seg_4_4_sp4_v_b_5_15247 = seg_3_4_sp4_r_v_b_5_15247;
  assign seg_4_4_sp4_v_b_6_15250 = net_15250;
  assign seg_4_4_sp4_v_b_7_15249 = seg_3_2_sp4_r_v_b_31_15249;
  assign seg_4_5_lutff_0_out_15593 = net_15593;
  assign seg_4_5_lutff_3_out_15596 = net_15596;
  assign seg_4_5_lutff_4_out_15597 = net_15597;
  assign seg_4_5_lutff_5_out_15598 = net_15598;
  assign seg_4_5_lutff_6_out_15599 = net_15599;
  assign seg_4_5_lutff_7_out_15600 = net_15600;
  assign seg_4_5_neigh_op_bnl_0_11639 = seg_3_4_lutff_0_out_11639;
  assign seg_4_5_neigh_op_bnr_6_19307 = seg_5_4_lutff_6_out_19307;
  assign seg_4_5_neigh_op_rgt_7_19431 = seg_5_5_lutff_7_out_19431;
  assign seg_4_5_sp4_h_l_37_1178 = seg_0_5_sp4_h_r_0_1178;
  assign seg_4_5_sp4_h_l_44_1225 = seg_1_5_sp4_h_r_20_1225;
  assign seg_4_5_sp4_h_r_10_19561 = net_19561;
  assign seg_4_5_sp4_h_r_12_15729 = net_15729;
  assign seg_4_5_sp4_h_r_18_15737 = net_15737;
  assign seg_4_5_sp4_h_r_20_15739 = net_15739;
  assign seg_4_5_sp4_h_r_28_11903 = net_11903;
  assign seg_4_5_sp4_v_b_28_15622 = net_15622;
  assign seg_4_5_sp4_v_b_42_15746 = net_15746;
  assign seg_4_5_sp4_v_b_44_15748 = net_15748;
  assign seg_4_6_lutff_0_out_15716 = net_15716;
  assign seg_4_6_lutff_1_out_15717 = net_15717;
  assign seg_4_6_lutff_2_out_15718 = net_15718;
  assign seg_4_6_lutff_3_out_15719 = net_15719;
  assign seg_4_6_lutff_5_out_15721 = net_15721;
  assign seg_4_6_lutff_6_out_15722 = net_15722;
  assign seg_4_6_lutff_7_out_15723 = net_15723;
  assign seg_4_6_neigh_op_lft_0_11885 = seg_3_6_lutff_0_out_11885;
  assign seg_4_6_sp4_h_l_37_1384 = seg_0_6_sp4_h_r_0_1384;
  assign seg_4_6_sp4_h_l_41_1418 = seg_0_6_sp4_h_r_4_1418;
  assign seg_4_6_sp4_h_l_47_1386 = seg_2_6_sp4_h_r_34_1386;
  assign seg_4_6_sp4_h_r_5_19689 = seg_7_6_sp4_h_r_40_19689;
  assign seg_4_6_sp4_h_r_9_19693 = seg_7_6_sp4_h_r_44_19693;
  assign seg_4_6_sp4_r_v_b_41_19699 = net_19699;
  assign seg_4_7_lutff_1_out_15840 = net_15840;
  assign seg_4_7_lutff_3_out_15842 = net_15842;
  assign seg_4_7_lutff_5_out_15844 = net_15844;
  assign seg_4_7_lutff_6_out_15845 = net_15845;
  assign seg_4_7_lutff_7_out_15846 = net_15846;
  assign seg_4_7_neigh_op_bnl_5_11890 = seg_3_6_lutff_5_out_11890;
  assign seg_4_7_neigh_op_bnl_7_11892 = seg_3_6_lutff_7_out_11892;
  assign seg_4_7_neigh_op_rgt_3_19673 = seg_5_7_lutff_3_out_19673;
  assign seg_4_7_sp4_h_l_43_1636 = seg_0_7_sp4_h_r_6_1636;
  assign seg_4_7_sp4_h_l_47_1594 = seg_0_7_sp4_h_r_10_1594;
  assign seg_4_7_sp4_h_r_0_19805 = net_19805;
  assign seg_4_7_sp4_h_r_4_19811 = net_19811;
  assign seg_4_7_sp4_r_v_b_9_19456 = net_19456;
  assign seg_4_7_sp4_v_b_18_15746 = seg_4_5_sp4_v_b_42_15746;
  assign seg_4_7_sp4_v_b_20_15748 = seg_4_5_sp4_v_b_44_15748;
  assign seg_4_7_sp4_v_t_36_16109 = seg_3_11_sp4_r_v_b_1_16109;
  assign seg_4_7_sp4_v_t_38_16111 = seg_3_11_sp4_r_v_b_3_16111;
  assign seg_4_7_sp4_v_t_42_16115 = seg_3_11_sp4_r_v_b_7_16115;
  assign seg_4_7_sp4_v_t_43_16116 = seg_4_11_sp4_v_b_6_16116;
  assign seg_4_7_sp4_v_t_45_16118 = seg_4_11_sp4_v_b_8_16118;
  assign seg_4_8_neigh_op_lft_4_12135 = seg_3_8_lutff_4_out_12135;
  assign seg_4_8_neigh_op_tnl_1_12255 = seg_3_9_lutff_1_out_12255;
  assign seg_4_8_neigh_op_tnl_2_12256 = seg_3_9_lutff_2_out_12256;
  assign seg_4_8_neigh_op_tnl_3_12257 = seg_3_9_lutff_3_out_12257;
  assign seg_4_8_neigh_op_tnl_4_12258 = seg_3_9_lutff_4_out_12258;
  assign seg_4_8_neigh_op_tnl_5_12259 = seg_3_9_lutff_5_out_12259;
  assign seg_4_8_neigh_op_tnl_6_12260 = seg_3_9_lutff_6_out_12260;
  assign seg_4_8_neigh_op_tnl_7_12261 = seg_3_9_lutff_7_out_12261;
  assign seg_4_8_sp12_h_r_1_19925 = seg_11_8_sp12_h_r_14_19925;
  assign seg_4_8_sp4_h_l_37_1801 = seg_0_8_sp4_h_r_0_1801;
  assign seg_4_8_sp4_r_v_b_47_19951 = net_19951;
  assign seg_4_8_sp4_v_t_40_16236 = seg_3_10_sp4_r_v_b_29_16236;
  assign seg_4_9_neigh_op_lft_7_12261 = seg_3_9_lutff_7_out_12261;
  assign seg_4_9_sp4_h_r_11_20054 = seg_5_9_sp4_h_r_22_20054;
  assign seg_4_9_sp4_h_r_14_16225 = net_16225;
  assign seg_4_9_sp4_h_r_20_16231 = net_16231;
  assign seg_4_9_sp4_h_r_22_16223 = net_16223;
  assign seg_4_9_sp4_h_r_24_12389 = net_12389;
  assign seg_4_9_sp4_h_r_32_12399 = net_12399;
  assign seg_4_9_sp4_h_r_5_20058 = seg_5_9_sp4_h_r_16_20058;
  assign seg_4_9_sp4_h_r_9_20062 = seg_5_9_sp4_h_r_20_20062;
  assign seg_4_9_sp4_r_v_b_27_19942 = net_19942;
  assign seg_4_9_sp4_r_v_b_29_19944 = net_19944;
  assign seg_4_9_sp4_r_v_b_35_19950 = net_19950;
  assign seg_4_9_sp4_v_t_45_16364 = seg_4_11_sp4_v_b_32_16364;
  assign seg_5_0_logic_op_top_7_18898 = seg_5_1_lutff_7_out_18898;
  assign seg_5_0_span4_horz_r_2_22756 = seg_6_0_span4_horz_r_6_22756;
  assign seg_5_10_sp12_v_b_12_23266 = net_23266;
  assign seg_5_10_sp12_v_b_4_22746 = seg_5_12_sp12_v_b_0_22746;
  assign seg_5_10_sp4_h_l_41_8202 = seg_1_10_sp4_h_r_4_8202;
  assign seg_5_10_sp4_h_r_10_24007 = net_24007;
  assign seg_5_10_sp4_h_r_16_20181 = net_20181;
  assign seg_5_10_sp4_h_r_1_24006 = seg_6_10_sp4_h_r_12_24006;
  assign seg_5_10_sp4_r_v_b_15_23774 = net_23774;
  assign seg_5_10_sp4_r_v_b_19_23778 = net_23778;
  assign seg_5_10_sp4_r_v_b_39_24020 = net_24020;
  assign seg_5_10_sp4_v_b_20_19948 = net_19948;
  assign seg_5_10_sp4_v_b_26_20066 = seg_5_12_sp4_v_b_2_20066;
  assign seg_5_10_sp4_v_b_40_20190 = net_20190;
  assign seg_5_10_sp4_v_t_39_20312 = seg_5_12_sp4_v_b_26_20312;
  assign seg_5_10_sp4_v_t_40_20313 = seg_5_13_sp4_v_b_16_20313;
  assign seg_5_10_sp4_v_t_44_20317 = seg_5_13_sp4_v_b_20_20317;
  assign seg_5_10_sp4_v_t_46_20319 = seg_5_11_sp4_v_b_46_20319;
  assign seg_5_11_neigh_op_rgt_0_23993 = seg_6_11_ram_RDATA_15_23993;
  assign seg_5_11_neigh_op_rgt_2_23995 = seg_6_11_ram_RDATA_13_23995;
  assign seg_5_11_neigh_op_rgt_4_23997 = seg_6_11_ram_RDATA_11_23997;
  assign seg_5_11_neigh_op_tnr_0_24116 = seg_6_12_ram_RDATA_7_24116;
  assign seg_5_11_neigh_op_tnr_4_24120 = seg_6_12_ram_RDATA_3_24120;
  assign seg_5_11_sp4_h_l_43_8351 = seg_1_11_sp4_h_r_6_8351;
  assign seg_5_11_sp4_h_r_18_20306 = net_20306;
  assign seg_5_11_sp4_h_r_32_16476 = net_16476;
  assign seg_5_11_sp4_h_r_6_24136 = net_24136;
  assign seg_5_11_sp4_r_v_b_10_23782 = seg_6_9_sp4_v_b_34_23782;
  assign seg_5_11_sp4_v_b_10_19951 = seg_4_8_sp4_r_v_b_47_19951;
  assign seg_5_11_sp4_v_b_11_19950 = seg_4_9_sp4_r_v_b_35_19950;
  assign seg_5_11_sp4_v_b_24_20187 = net_20187;
  assign seg_5_11_sp4_v_b_26_20189 = net_20189;
  assign seg_5_11_sp4_v_b_28_20191 = net_20191;
  assign seg_5_11_sp4_v_b_32_20195 = net_20195;
  assign seg_5_11_sp4_v_b_36_20309 = net_20309;
  assign seg_5_11_sp4_v_b_3_19942 = seg_4_9_sp4_r_v_b_27_19942;
  assign seg_5_11_sp4_v_b_46_20319 = net_20319;
  assign seg_5_11_sp4_v_b_4_19945 = net_19945;
  assign seg_5_11_sp4_v_b_5_19944 = seg_4_9_sp4_r_v_b_29_19944;
  assign seg_5_11_sp4_v_b_9_19948 = seg_5_10_sp4_v_b_20_19948;
  assign seg_5_12_lutff_2_out_20287 = net_20287;
  assign seg_5_12_lutff_4_out_20289 = net_20289;
  assign seg_5_12_neigh_op_bnr_5_23998 = seg_6_11_ram_RDATA_10_23998;
  assign seg_5_12_neigh_op_top_4_20412 = seg_5_13_lutff_4_out_20412;
  assign seg_5_12_neigh_op_top_7_20415 = seg_5_13_lutff_7_out_20415;
  assign seg_5_12_sp12_v_b_0_22746 = net_22746;
  assign seg_5_12_sp4_h_r_18_20429 = net_20429;
  assign seg_5_12_sp4_h_r_22_20423 = net_20423;
  assign seg_5_12_sp4_h_r_28_16595 = net_16595;
  assign seg_5_12_sp4_h_r_32_16599 = net_16599;
  assign seg_5_12_sp4_h_r_34_16591 = net_16591;
  assign seg_5_12_sp4_h_r_3_24256 = seg_6_12_sp4_h_r_14_24256;
  assign seg_5_12_sp4_h_r_46_12761 = net_12761;
  assign seg_5_12_sp4_r_v_b_19_24024 = net_24024;
  assign seg_5_12_sp4_r_v_b_31_24146 = net_24146;
  assign seg_5_12_sp4_r_v_b_33_24148 = net_24148;
  assign seg_5_12_sp4_v_b_11_20073 = seg_5_9_sp4_v_b_46_20073;
  assign seg_5_12_sp4_v_b_1_20063 = seg_5_9_sp4_v_b_36_20063;
  assign seg_5_12_sp4_v_b_26_20312 = net_20312;
  assign seg_5_12_sp4_v_b_2_20066 = net_20066;
  assign seg_5_12_sp4_v_b_3_20065 = seg_5_9_sp4_v_b_38_20065;
  assign seg_5_12_sp4_v_b_41_20437 = seg_5_15_sp4_v_b_4_20437;
  assign seg_5_12_sp4_v_b_5_20067 = seg_5_9_sp4_v_b_40_20067;
  assign seg_5_12_sp4_v_b_6_20070 = net_20070;
  assign seg_5_12_sp4_v_b_7_20069 = seg_5_9_sp4_v_b_42_20069;
  assign seg_5_12_sp4_v_b_9_20071 = seg_5_9_sp4_v_b_44_20071;
  assign seg_5_12_sp4_v_t_41_20560 = seg_5_16_sp4_v_b_4_20560;
  assign seg_5_12_sp4_v_t_47_20566 = seg_5_16_sp4_v_b_10_20566;
  assign seg_5_13_lutff_0_out_20408 = net_20408;
  assign seg_5_13_lutff_2_out_20410 = net_20410;
  assign seg_5_13_lutff_3_out_20411 = net_20411;
  assign seg_5_13_lutff_4_out_20412 = net_20412;
  assign seg_5_13_lutff_5_out_20413 = net_20413;
  assign seg_5_13_lutff_6_out_20414 = net_20414;
  assign seg_5_13_lutff_7_out_20415 = net_20415;
  assign seg_5_13_sp12_v_b_0_22861 = net_22861;
  assign seg_5_13_sp4_h_r_18_20552 = net_20552;
  assign seg_5_13_sp4_h_r_26_16716 = seg_3_13_sp4_h_r_2_16716;
  assign seg_5_13_sp4_h_r_32_16722 = seg_3_13_sp4_h_r_8_16722;
  assign seg_5_13_sp4_h_r_34_16714 = seg_3_13_sp4_h_r_10_16714;
  assign seg_5_13_sp4_h_r_44_12892 = seg_3_13_sp4_h_r_20_12892;
  assign seg_5_13_sp4_h_r_46_12884 = seg_3_13_sp4_h_r_22_12884;
  assign seg_5_13_sp4_r_v_b_17_24145 = net_24145;
  assign seg_5_13_sp4_r_v_b_19_24147 = net_24147;
  assign seg_5_13_sp4_v_b_0_20187 = seg_5_11_sp4_v_b_24_20187;
  assign seg_5_13_sp4_v_b_10_20197 = seg_4_10_sp4_r_v_b_47_20197;
  assign seg_5_13_sp4_v_b_16_20313 = net_20313;
  assign seg_5_13_sp4_v_b_1_20186 = seg_4_11_sp4_r_v_b_25_20186;
  assign seg_5_13_sp4_v_b_20_20317 = net_20317;
  assign seg_5_13_sp4_v_b_2_20189 = seg_5_11_sp4_v_b_26_20189;
  assign seg_5_13_sp4_v_b_34_20443 = net_20443;
  assign seg_5_13_sp4_v_b_4_20191 = seg_5_11_sp4_v_b_28_20191;
  assign seg_5_13_sp4_v_b_5_20190 = seg_5_10_sp4_v_b_40_20190;
  assign seg_5_13_sp4_v_b_8_20195 = seg_5_11_sp4_v_b_32_20195;
  assign seg_5_14_lutff_1_out_20532 = net_20532;
  assign seg_5_14_lutff_2_out_20533 = net_20533;
  assign seg_5_14_lutff_4_out_20535 = net_20535;
  assign seg_5_14_lutff_5_out_20536 = net_20536;
  assign seg_5_14_sp4_h_l_36_8785 = seg_2_14_sp4_h_r_12_8785;
  assign seg_5_14_sp4_r_v_b_17_24268 = net_24268;
  assign seg_5_14_sp4_r_v_b_31_24392 = net_24392;
  assign seg_5_14_sp4_v_b_11_20319 = seg_5_11_sp4_v_b_46_20319;
  assign seg_5_14_sp4_v_b_1_20309 = seg_5_11_sp4_v_b_36_20309;
  assign seg_5_14_sp4_v_b_2_20312 = seg_5_12_sp4_v_b_26_20312;
  assign seg_5_14_sp4_v_t_41_20806 = seg_5_16_sp4_v_b_28_20806;
  assign seg_5_15_lutff_1_out_20655 = net_20655;
  assign seg_5_15_lutff_3_out_20657 = net_20657;
  assign seg_5_15_lutff_4_out_20658 = net_20658;
  assign seg_5_15_lutff_6_out_20660 = net_20660;
  assign seg_5_15_lutff_7_out_20661 = net_20661;
  assign seg_5_15_sp4_r_v_b_43_24639 = net_24639;
  assign seg_5_15_sp4_v_b_10_20443 = seg_5_13_sp4_v_b_34_20443;
  assign seg_5_15_sp4_v_b_2_20435 = seg_4_12_sp4_r_v_b_39_20435;
  assign seg_5_15_sp4_v_b_4_20437 = net_20437;
  assign seg_5_15_sp4_v_t_42_20930 = seg_4_17_sp4_r_v_b_31_20930;
  assign seg_5_16_sp12_v_b_0_23266 = seg_5_10_sp12_v_b_12_23266;
  assign seg_5_16_sp12_v_b_3_23389 = seg_5_7_sp12_v_b_20_23389;
  assign seg_5_16_sp4_r_v_b_15_24512 = net_24512;
  assign seg_5_16_sp4_r_v_b_27_24634 = seg_5_18_sp4_r_v_b_3_24634;
  assign seg_5_16_sp4_v_b_10_20566 = net_20566;
  assign seg_5_16_sp4_v_b_28_20806 = net_20806;
  assign seg_5_16_sp4_v_b_4_20560 = net_20560;
  assign seg_5_17_lutff_1_out_20901 = net_20901;
  assign seg_5_17_sp4_h_r_2_24870 = net_24870;
  assign seg_5_17_sp4_h_r_34_17206 = net_17206;
  assign seg_5_18_neigh_op_tnl_6_17321 = seg_4_19_lutff_6_out_17321;
  assign seg_5_18_neigh_op_top_0_21146 = seg_5_19_lutff_0_out_21146;
  assign seg_5_18_sp4_h_r_22_21161 = net_21161;
  assign seg_5_18_sp4_h_r_24_17327 = net_17327;
  assign seg_5_18_sp4_r_v_b_3_24634 = net_24634;
  assign seg_5_19_lutff_0_out_21146 = net_21146;
  assign seg_5_19_neigh_op_tnl_4_17442 = seg_4_20_lutff_4_out_17442;
  assign seg_5_19_sp12_v_t_23_25111 = seg_5_31_span12_vert_0_25111;
  assign seg_5_19_sp4_h_r_24_17450 = net_17450;
  assign seg_5_1_lutff_3_out_18894 = net_18894;
  assign seg_5_1_lutff_7_out_18898 = net_18898;
  assign seg_5_1_sp4_v_b_42_19080 = seg_4_4_sp4_r_v_b_7_19080;
  assign seg_5_2_lutff_5_out_19024 = net_19024;
  assign seg_5_2_sp12_v_b_20_22746 = seg_5_12_sp12_v_b_0_22746;
  assign seg_5_2_sp4_h_l_46_7023 = seg_2_2_sp4_h_r_22_7023;
  assign seg_5_2_sp4_r_v_b_19_22898 = net_22898;
  assign seg_5_30_sp4_v_t_40_26489 = seg_5_31_span4_vert_40_26489;
  assign seg_5_31_span12_vert_0_25111 = net_25111;
  assign seg_5_31_span4_vert_40_26489 = net_26489;
  assign seg_5_3_lutff_2_out_19180 = net_19180;
  assign seg_5_3_lutff_5_out_19183 = net_19183;
  assign seg_5_3_neigh_op_bot_5_19024 = seg_5_2_lutff_5_out_19024;
  assign seg_5_3_sp12_v_b_19_22746 = seg_5_12_sp12_v_b_0_22746;
  assign seg_5_3_sp12_v_b_20_22861 = seg_5_13_sp12_v_b_0_22861;
  assign seg_5_3_sp4_h_l_42_7176 = seg_4_3_sp4_h_r_42_7176;
  assign seg_5_3_sp4_h_l_45_7177 = seg_1_3_sp4_h_r_8_7177;
  assign seg_5_3_sp4_h_l_47_7169 = seg_1_3_sp4_h_r_10_7169;
  assign seg_5_3_sp4_v_b_30_19209 = net_19209;
  assign seg_5_3_sp4_v_b_8_19069 = net_19069;
  assign seg_5_3_sp4_v_t_44_19456 = seg_4_7_sp4_r_v_b_9_19456;
  assign seg_5_4_lutff_6_out_19307 = net_19307;
  assign seg_5_4_neigh_op_bnr_4_23013 = seg_6_3_ram_RDATA_11_23013;
  assign seg_5_4_neigh_op_bnr_5_23014 = seg_6_3_ram_RDATA_10_23014;
  assign seg_5_4_neigh_op_bnr_6_23015 = seg_6_3_ram_RDATA_9_23015;
  assign seg_5_4_neigh_op_bnr_7_23016 = seg_6_3_ram_RDATA_8_23016;
  assign seg_5_4_neigh_op_rgt_0_23132 = seg_6_4_ram_RDATA_7_23132;
  assign seg_5_4_neigh_op_rgt_1_23133 = seg_6_4_ram_RDATA_6_23133;
  assign seg_5_4_neigh_op_tnl_7_15600 = seg_4_5_lutff_7_out_15600;
  assign seg_5_4_sp4_h_r_14_19441 = net_19441;
  assign seg_5_4_sp4_h_r_4_23273 = net_23273;
  assign seg_5_4_sp4_r_v_b_43_23286 = net_23286;
  assign seg_5_4_sp4_r_v_b_45_23288 = net_23288;
  assign seg_5_4_sp4_v_b_24_19326 = net_19326;
  assign seg_5_4_sp4_v_b_32_19334 = net_19334;
  assign seg_5_4_sp4_v_b_34_19336 = net_19336;
  assign seg_5_4_sp4_v_b_36_19448 = net_19448;
  assign seg_5_4_sp4_v_b_38_19450 = net_19450;
  assign seg_5_4_sp4_v_b_6_19081 = seg_4_1_sp4_r_v_b_43_19081;
  assign seg_5_5_lutff_7_out_19431 = net_19431;
  assign seg_5_5_neigh_op_lft_3_15596 = seg_4_5_lutff_3_out_15596;
  assign seg_5_5_neigh_op_top_1_19548 = seg_5_6_lutff_1_out_19548;
  assign seg_5_5_neigh_op_top_2_19549 = seg_5_6_lutff_2_out_19549;
  assign seg_5_5_neigh_op_top_3_19550 = seg_5_6_lutff_3_out_19550;
  assign seg_5_5_neigh_op_top_4_19551 = seg_5_6_lutff_4_out_19551;
  assign seg_5_5_neigh_op_top_5_19552 = seg_5_6_lutff_5_out_19552;
  assign seg_5_5_neigh_op_top_6_19553 = seg_5_6_lutff_6_out_19553;
  assign seg_5_5_sp4_h_l_39_7465 = seg_3_5_sp4_h_r_26_7465;
  assign seg_5_5_sp4_h_r_0_23390 = seg_7_5_sp4_h_r_24_23390;
  assign seg_5_5_sp4_h_r_10_23392 = net_23392;
  assign seg_5_5_sp4_h_r_1_23391 = seg_8_5_sp4_h_r_36_23391;
  assign seg_5_5_sp4_h_r_34_15730 = net_15730;
  assign seg_5_5_sp4_h_r_36_11898 = net_11898;
  assign seg_5_5_sp4_h_r_38_11902 = net_11902;
  assign seg_5_5_sp4_h_r_40_11904 = net_11904;
  assign seg_5_5_sp4_r_v_b_13_23157 = net_23157;
  assign seg_5_5_sp4_v_b_6_19209 = seg_5_3_sp4_v_b_30_19209;
  assign seg_5_6_lutff_1_out_19548 = net_19548;
  assign seg_5_6_lutff_2_out_19549 = net_19549;
  assign seg_5_6_lutff_3_out_19550 = net_19550;
  assign seg_5_6_lutff_4_out_19551 = net_19551;
  assign seg_5_6_lutff_5_out_19552 = net_19552;
  assign seg_5_6_lutff_6_out_19553 = net_19553;
  assign seg_5_6_neigh_op_bnl_0_15593 = seg_4_5_lutff_0_out_15593;
  assign seg_5_6_sp4_h_r_10_23515 = seg_7_6_sp4_h_r_34_23515;
  assign seg_5_6_sp4_h_r_2_23517 = seg_7_6_sp4_h_r_26_23517;
  assign seg_5_6_sp4_h_r_30_15859 = net_15859;
  assign seg_5_6_sp4_r_v_b_19_23286 = seg_5_4_sp4_r_v_b_43_23286;
  assign seg_5_6_sp4_r_v_b_21_23288 = seg_5_4_sp4_r_v_b_45_23288;
  assign seg_5_6_sp4_v_b_0_19326 = seg_5_4_sp4_v_b_24_19326;
  assign seg_5_6_sp4_v_b_10_19336 = seg_5_4_sp4_v_b_34_19336;
  assign seg_5_6_sp4_v_b_12_19448 = seg_5_4_sp4_v_b_36_19448;
  assign seg_5_6_sp4_v_b_14_19450 = seg_5_4_sp4_v_b_38_19450;
  assign seg_5_6_sp4_v_b_26_19574 = seg_5_8_sp4_v_b_2_19574;
  assign seg_5_6_sp4_v_b_8_19334 = seg_5_4_sp4_v_b_32_19334;
  assign seg_5_7_lutff_3_out_19673 = net_19673;
  assign seg_5_7_neigh_op_lft_1_15840 = seg_4_7_lutff_1_out_15840;
  assign seg_5_7_neigh_op_lft_5_15844 = seg_4_7_lutff_5_out_15844;
  assign seg_5_7_neigh_op_top_3_19796 = seg_5_8_lutff_3_out_19796;
  assign seg_5_7_sp12_v_b_20_23389 = net_23389;
  assign seg_5_7_sp4_h_r_0_23636 = seg_7_7_sp4_h_r_24_23636;
  assign seg_5_7_sp4_h_r_18_19814 = net_19814;
  assign seg_5_7_sp4_h_r_2_23640 = seg_7_7_sp4_h_r_26_23640;
  assign seg_5_7_sp4_r_v_b_11_23289 = net_23289;
  assign seg_5_7_sp4_v_t_41_19945 = seg_5_11_sp4_v_b_4_19945;
  assign seg_5_8_lutff_3_out_19796 = net_19796;
  assign seg_5_8_lutff_5_out_19798 = net_19798;
  assign seg_5_8_lutff_6_out_19799 = net_19799;
  assign seg_5_8_neigh_op_bnl_3_15842 = seg_4_7_lutff_3_out_15842;
  assign seg_5_8_neigh_op_bot_3_19673 = seg_5_7_lutff_3_out_19673;
  assign seg_5_8_sp4_h_l_47_7904 = seg_1_8_sp4_h_r_10_7904;
  assign seg_5_8_sp4_h_r_14_19933 = net_19933;
  assign seg_5_8_sp4_h_r_20_19939 = net_19939;
  assign seg_5_8_sp4_h_r_6_23767 = net_23767;
  assign seg_5_8_sp4_h_r_8_23769 = net_23769;
  assign seg_5_8_sp4_r_v_b_1_23402 = net_23402;
  assign seg_5_8_sp4_r_v_b_23_23536 = net_23536;
  assign seg_5_8_sp4_v_b_2_19574 = net_19574;
  assign seg_5_8_sp4_v_t_39_20066 = seg_5_12_sp4_v_b_2_20066;
  assign seg_5_8_sp4_v_t_43_20070 = seg_5_12_sp4_v_b_6_20070;
  assign seg_5_8_sp4_v_t_46_20073 = seg_5_9_sp4_v_b_46_20073;
  assign seg_5_9_neigh_op_rgt_0_23747 = seg_6_9_ram_RDATA_15_23747;
  assign seg_5_9_neigh_op_rgt_2_23749 = seg_6_9_ram_RDATA_13_23749;
  assign seg_5_9_neigh_op_rgt_5_23752 = seg_6_9_ram_RDATA_10_23752;
  assign seg_5_9_neigh_op_tnr_0_23870 = seg_6_10_ram_RDATA_7_23870;
  assign seg_5_9_neigh_op_tnr_1_23871 = seg_6_10_ram_RDATA_6_23871;
  assign seg_5_9_neigh_op_tnr_2_23872 = seg_6_10_ram_RDATA_5_23872;
  assign seg_5_9_neigh_op_tnr_3_23873 = seg_6_10_ram_RDATA_4_23873;
  assign seg_5_9_neigh_op_tnr_7_23877 = seg_6_10_ram_RDATA_0_23877;
  assign seg_5_9_sp12_h_r_10_1991 = net_1991;
  assign seg_5_9_sp4_h_l_36_8050 = seg_2_9_sp4_h_r_12_8050;
  assign seg_5_9_sp4_h_l_46_8052 = seg_2_9_sp4_h_r_22_8052;
  assign seg_5_9_sp4_h_r_0_23882 = seg_7_9_sp4_h_r_24_23882;
  assign seg_5_9_sp4_h_r_16_20058 = net_20058;
  assign seg_5_9_sp4_h_r_20_20062 = net_20062;
  assign seg_5_9_sp4_h_r_22_20054 = net_20054;
  assign seg_5_9_sp4_r_v_b_25_23771 = net_23771;
  assign seg_5_9_sp4_r_v_b_27_23773 = net_23773;
  assign seg_5_9_sp4_r_v_b_29_23775 = net_23775;
  assign seg_5_9_sp4_r_v_b_33_23779 = net_23779;
  assign seg_5_9_sp4_r_v_b_35_23781 = net_23781;
  assign seg_5_9_sp4_v_b_36_20063 = net_20063;
  assign seg_5_9_sp4_v_b_38_20065 = net_20065;
  assign seg_5_9_sp4_v_b_40_20067 = net_20067;
  assign seg_5_9_sp4_v_b_42_20069 = net_20069;
  assign seg_5_9_sp4_v_b_44_20071 = net_20071;
  assign seg_5_9_sp4_v_b_46_20073 = net_20073;
  assign seg_5_9_sp4_v_b_4_19699 = seg_4_6_sp4_r_v_b_41_19699;
  assign seg_5_9_sp4_v_t_37_20187 = seg_5_11_sp4_v_b_24_20187;
  assign seg_5_9_sp4_v_t_39_20189 = seg_5_11_sp4_v_b_26_20189;
  assign seg_5_9_sp4_v_t_41_20191 = seg_5_11_sp4_v_b_28_20191;
  assign seg_6_0_span4_horz_r_6_22756 = net_22756;
  assign seg_6_0_span4_horz_r_8_18923 = net_18923;
  assign seg_6_0_span4_vert_0_22874 = net_22874;
  assign seg_6_0_span4_vert_28_22895 = net_22895;
  assign seg_6_10_ram_RDATA_0_23877 = net_23877;
  assign seg_6_10_ram_RDATA_4_23873 = net_23873;
  assign seg_6_10_ram_RDATA_5_23872 = net_23872;
  assign seg_6_10_ram_RDATA_6_23871 = net_23871;
  assign seg_6_10_ram_RDATA_7_23870 = net_23870;
  assign seg_6_10_sp4_h_r_10_27627 = net_27627;
  assign seg_6_10_sp4_h_r_12_24006 = net_24006;
  assign seg_6_10_sp4_h_r_8_27635 = net_27635;
  assign seg_6_10_sp4_v_t_41_24145 = seg_5_13_sp4_r_v_b_17_24145;
  assign seg_6_10_sp4_v_t_42_24146 = seg_5_12_sp4_r_v_b_31_24146;
  assign seg_6_10_sp4_v_t_43_24147 = seg_5_13_sp4_r_v_b_19_24147;
  assign seg_6_10_sp4_v_t_44_24148 = seg_5_12_sp4_r_v_b_33_24148;
  assign seg_6_11_ram_RDATA_10_23998 = net_23998;
  assign seg_6_11_ram_RDATA_11_23997 = net_23997;
  assign seg_6_11_ram_RDATA_13_23995 = net_23995;
  assign seg_6_11_ram_RDATA_15_23993 = net_23993;
  assign seg_6_11_sp4_h_r_2_27731 = net_27731;
  assign seg_6_11_sp4_h_r_38_16471 = net_16471;
  assign seg_6_11_sp4_h_r_44_16477 = net_16477;
  assign seg_6_11_sp4_h_r_46_16469 = net_16469;
  assign seg_6_11_sp4_h_r_9_27738 = seg_9_11_sp4_h_r_44_27738;
  assign seg_6_11_sp4_v_b_11_23781 = seg_5_9_sp4_r_v_b_35_23781;
  assign seg_6_11_sp4_v_b_1_23771 = seg_5_9_sp4_r_v_b_25_23771;
  assign seg_6_11_sp4_v_b_2_23774 = seg_5_10_sp4_r_v_b_15_23774;
  assign seg_6_11_sp4_v_b_3_23773 = seg_5_9_sp4_r_v_b_27_23773;
  assign seg_6_11_sp4_v_b_5_23775 = seg_5_9_sp4_r_v_b_29_23775;
  assign seg_6_11_sp4_v_b_6_23778 = seg_5_10_sp4_r_v_b_19_23778;
  assign seg_6_11_sp4_v_b_9_23779 = seg_5_9_sp4_r_v_b_33_23779;
  assign seg_6_11_sp4_v_t_36_24263 = seg_6_12_sp4_v_b_36_24263;
  assign seg_6_11_sp4_v_t_38_24265 = seg_6_12_sp4_v_b_38_24265;
  assign seg_6_11_sp4_v_t_41_24268 = seg_5_14_sp4_r_v_b_17_24268;
  assign seg_6_12_ram_RDATA_3_24120 = net_24120;
  assign seg_6_12_ram_RDATA_7_24116 = net_24116;
  assign seg_6_12_sp4_h_r_14_24256 = net_24256;
  assign seg_6_12_sp4_h_r_28_20426 = net_20426;
  assign seg_6_12_sp4_h_r_34_20422 = net_20422;
  assign seg_6_12_sp4_v_b_10_23905 = net_23905;
  assign seg_6_12_sp4_v_b_36_24263 = net_24263;
  assign seg_6_12_sp4_v_b_38_24265 = net_24265;
  assign seg_6_12_sp4_v_t_42_24392 = seg_5_14_sp4_r_v_b_31_24392;
  assign seg_6_13_sp4_h_l_36_12882 = seg_3_13_sp4_h_r_12_12882;
  assign seg_6_13_sp4_h_l_47_12883 = seg_2_13_sp4_h_r_10_12883;
  assign seg_6_13_sp4_v_b_2_24020 = seg_5_10_sp4_r_v_b_39_24020;
  assign seg_6_13_sp4_v_t_39_24512 = seg_5_16_sp4_r_v_b_15_24512;
  assign seg_6_14_sp4_v_t_43_24639 = seg_5_15_sp4_r_v_b_43_24639;
  assign seg_6_19_sp12_v_t_23_28542 = seg_6_31_span12_vert_0_28542;
  assign seg_6_1_sp4_h_l_36_11370 = seg_3_1_sp4_h_r_12_11370;
  assign seg_6_1_sp4_h_l_38_11374 = seg_3_1_sp4_h_r_14_11374;
  assign seg_6_1_sp4_h_l_42_11378 = seg_3_1_sp4_h_r_18_11378;
  assign seg_6_1_sp4_h_l_44_11380 = seg_3_1_sp4_h_r_20_11380;
  assign seg_6_1_sp4_v_b_0_22874 = seg_6_0_span4_vert_0_22874;
  assign seg_6_28_sp4_v_t_40_26358 = seg_6_31_span4_vert_16_26358;
  assign seg_6_2_sp4_h_l_37_11528 = seg_2_2_sp4_h_r_0_11528;
  assign seg_6_2_sp4_h_l_43_11536 = seg_2_2_sp4_h_r_6_11536;
  assign seg_6_2_sp4_h_l_45_11538 = seg_2_2_sp4_h_r_8_11538;
  assign seg_6_30_sp4_v_t_40_29689 = seg_6_31_span4_vert_40_29689;
  assign seg_6_31_span12_vert_0_28542 = net_28542;
  assign seg_6_31_span4_vert_16_26358 = net_26358;
  assign seg_6_31_span4_vert_40_29689 = net_29689;
  assign seg_6_3_neigh_op_lft_2_19180 = seg_5_3_lutff_2_out_19180;
  assign seg_6_3_ram_RDATA_10_23014 = net_23014;
  assign seg_6_3_ram_RDATA_11_23013 = net_23013;
  assign seg_6_3_ram_RDATA_8_23016 = net_23016;
  assign seg_6_3_ram_RDATA_9_23015 = net_23015;
  assign seg_6_3_sp4_h_r_41_15488 = seg_3_3_sp4_h_r_4_15488;
  assign seg_6_3_sp4_h_r_43_15490 = seg_3_3_sp4_h_r_6_15490;
  assign seg_6_3_sp4_v_b_4_22895 = seg_6_0_span4_vert_28_22895;
  assign seg_6_3_sp4_v_b_6_22898 = seg_5_2_sp4_r_v_b_19_22898;
  assign seg_6_4_neigh_op_bnl_2_19180 = seg_5_3_lutff_2_out_19180;
  assign seg_6_4_ram_RDATA_6_23133 = net_23133;
  assign seg_6_4_ram_RDATA_7_23132 = net_23132;
  assign seg_6_4_sp4_h_l_36_11775 = seg_3_4_sp4_h_r_12_11775;
  assign seg_6_4_sp4_h_l_39_11778 = seg_4_4_sp4_h_r_26_11778;
  assign seg_6_4_sp4_h_l_47_11776 = seg_2_4_sp4_h_r_10_11776;
  assign seg_6_4_sp4_h_r_36_15606 = net_15606;
  assign seg_6_4_sp4_h_r_46_15608 = net_15608;
  assign seg_6_4_sp4_r_v_b_39_27028 = net_27028;
  assign seg_6_4_sp4_r_v_b_43_27032 = net_27032;
  assign seg_6_4_sp4_v_b_40_23283 = net_23283;
  assign seg_6_4_sp4_v_b_44_23287 = net_23287;
  assign seg_6_4_sp4_v_t_36_23402 = seg_5_8_sp4_r_v_b_1_23402;
  assign seg_6_5_sp4_h_l_41_11903 = seg_4_5_sp4_h_r_28_11903;
  assign seg_6_5_sp4_v_t_47_23536 = seg_5_8_sp4_r_v_b_23_23536;
  assign seg_6_6_sp4_h_l_36_12021 = seg_3_6_sp4_h_r_12_12021;
  assign seg_6_6_sp4_h_l_47_12022 = seg_2_6_sp4_h_r_10_12022;
  assign seg_6_6_sp4_v_b_0_23157 = seg_5_5_sp4_r_v_b_13_23157;
  assign seg_6_7_sp4_v_b_11_23289 = seg_5_7_sp4_r_v_b_11_23289;
  assign seg_6_7_sp4_v_b_5_23283 = seg_6_4_sp4_v_b_40_23283;
  assign seg_6_7_sp4_v_b_9_23287 = seg_6_4_sp4_v_b_44_23287;
  assign seg_6_8_sp4_h_l_43_12274 = seg_2_8_sp4_h_r_6_12274;
  assign seg_6_8_sp4_h_l_44_12277 = seg_3_8_sp4_h_r_20_12277;
  assign seg_6_8_sp4_h_l_45_12276 = seg_2_8_sp4_h_r_8_12276;
  assign seg_6_9_ram_RDATA_10_23752 = net_23752;
  assign seg_6_9_ram_RDATA_13_23749 = net_23749;
  assign seg_6_9_ram_RDATA_15_23747 = net_23747;
  assign seg_6_9_sp12_h_r_14_2002 = net_2002;
  assign seg_6_9_sp12_h_r_20_2012 = net_2012;
  assign seg_6_9_sp12_h_r_22_1992 = net_1992;
  assign seg_6_9_sp4_h_r_1_27524 = seg_7_9_sp4_h_r_12_27524;
  assign seg_6_9_sp4_h_r_40_16227 = net_16227;
  assign seg_6_9_sp4_v_b_34_23782 = net_23782;
  assign seg_6_9_sp4_v_t_43_24024 = seg_5_12_sp4_r_v_b_19_24024;
  assign seg_7_10_lutff_0_out_27481 = net_27481;
  assign seg_7_10_lutff_1_out_27482 = net_27482;
  assign seg_7_10_lutff_2_out_27483 = net_27483;
  assign seg_7_10_lutff_4_out_27485 = net_27485;
  assign seg_7_10_lutff_6_out_27487 = net_27487;
  assign seg_7_10_sp4_h_l_41_16349 = seg_3_10_sp4_h_r_4_16349;
  assign seg_7_10_sp4_v_b_46_27647 = net_27647;
  assign seg_7_10_sp4_v_b_6_27338 = net_27338;
  assign seg_7_10_sp4_v_t_36_27739 = seg_7_13_sp4_v_b_12_27739;
  assign seg_7_10_sp4_v_t_43_27746 = seg_7_14_sp4_v_b_6_27746;
  assign seg_7_11_lutff_0_out_27583 = net_27583;
  assign seg_7_11_lutff_1_out_27584 = net_27584;
  assign seg_7_11_lutff_2_out_27585 = net_27585;
  assign seg_7_11_lutff_3_out_27586 = net_27586;
  assign seg_7_11_lutff_6_out_27589 = net_27589;
  assign seg_7_11_lutff_7_out_27590 = net_27590;
  assign seg_7_11_neigh_op_bot_6_27487 = seg_7_10_lutff_6_out_27487;
  assign seg_7_11_sp4_h_r_30_24136 = seg_5_11_sp4_h_r_6_24136;
  assign seg_7_11_sp4_h_r_42_20306 = seg_5_11_sp4_h_r_18_20306;
  assign seg_7_11_sp4_h_r_4_31165 = seg_9_11_sp4_h_r_28_31165;
  assign seg_7_11_sp4_h_r_8_31169 = seg_9_11_sp4_h_r_32_31169;
  assign seg_7_11_sp4_v_b_10_27444 = seg_7_9_sp4_v_b_34_27444;
  assign seg_7_11_sp4_v_b_26_27640 = net_27640;
  assign seg_7_11_sp4_v_b_3_27435 = seg_7_8_sp4_v_b_38_27435;
  assign seg_7_11_sp4_v_b_40_27743 = net_27743;
  assign seg_7_11_sp4_v_t_39_27844 = seg_7_15_sp4_v_b_2_27844;
  assign seg_7_11_sp4_v_t_45_27850 = seg_7_15_sp4_v_b_8_27850;
  assign seg_7_12_lutff_1_out_27686 = net_27686;
  assign seg_7_12_lutff_2_out_27687 = net_27687;
  assign seg_7_12_lutff_3_out_27688 = net_27688;
  assign seg_7_12_lutff_4_out_27689 = net_27689;
  assign seg_7_12_lutff_5_out_27690 = net_27690;
  assign seg_7_12_lutff_6_out_27691 = net_27691;
  assign seg_7_12_lutff_7_out_27692 = net_27692;
  assign seg_7_12_neigh_op_bnr_1_31025 = seg_8_11_lutff_1_out_31025;
  assign seg_7_12_neigh_op_bnr_3_31027 = seg_8_11_lutff_3_out_31027;
  assign seg_7_12_neigh_op_bot_0_27583 = seg_7_11_lutff_0_out_27583;
  assign seg_7_12_neigh_op_bot_1_27584 = seg_7_11_lutff_1_out_27584;
  assign seg_7_12_neigh_op_bot_2_27585 = seg_7_11_lutff_2_out_27585;
  assign seg_7_12_neigh_op_bot_3_27586 = seg_7_11_lutff_3_out_27586;
  assign seg_7_12_neigh_op_bot_7_27590 = seg_7_11_lutff_7_out_27590;
  assign seg_7_12_neigh_op_tnr_3_31273 = seg_8_13_lutff_3_out_31273;
  assign seg_7_12_neigh_op_tnr_5_31275 = seg_8_13_lutff_5_out_31275;
  assign seg_7_12_neigh_op_top_2_27789 = seg_7_13_lutff_2_out_27789;
  assign seg_7_12_neigh_op_top_4_27791 = seg_7_13_lutff_4_out_27791;
  assign seg_7_12_neigh_op_top_5_27792 = seg_7_13_lutff_5_out_27792;
  assign seg_7_12_neigh_op_top_7_27794 = seg_7_13_lutff_7_out_27794;
  assign seg_7_12_sp4_h_l_42_16598 = seg_4_12_sp4_h_r_18_16598;
  assign seg_7_12_sp4_h_l_45_16599 = seg_5_12_sp4_h_r_32_16599;
  assign seg_7_12_sp4_r_v_b_18_31054 = seg_7_13_sp4_r_v_b_7_31054;
  assign seg_7_12_sp4_v_b_1_27535 = seg_7_9_sp4_v_b_36_27535;
  assign seg_7_12_sp4_v_b_3_27537 = seg_7_9_sp4_v_b_38_27537;
  assign seg_7_12_sp4_v_t_36_27943 = seg_7_15_sp4_v_b_12_27943;
  assign seg_7_13_lutff_0_out_27787 = net_27787;
  assign seg_7_13_lutff_1_out_27788 = net_27788;
  assign seg_7_13_lutff_2_out_27789 = net_27789;
  assign seg_7_13_lutff_4_out_27791 = net_27791;
  assign seg_7_13_lutff_5_out_27792 = net_27792;
  assign seg_7_13_lutff_7_out_27794 = net_27794;
  assign seg_7_13_sp4_h_l_38_16717 = seg_4_13_sp4_h_r_14_16717;
  assign seg_7_13_sp4_r_v_b_13_31172 = net_31172;
  assign seg_7_13_sp4_r_v_b_7_31054 = net_31054;
  assign seg_7_13_sp4_v_b_11_27647 = seg_7_10_sp4_v_b_46_27647;
  assign seg_7_13_sp4_v_b_12_27739 = net_27739;
  assign seg_7_13_sp4_v_b_16_27743 = seg_7_11_sp4_v_b_40_27743;
  assign seg_7_13_sp4_v_b_2_27640 = seg_7_11_sp4_v_b_26_27640;
  assign seg_7_14_lutff_6_out_27895 = net_27895;
  assign seg_7_14_lutff_7_out_27896 = net_27896;
  assign seg_7_14_neigh_op_top_2_27993 = seg_7_15_lutff_2_out_27993;
  assign seg_7_14_sp4_h_r_22_28036 = net_28036;
  assign seg_7_14_sp4_r_v_b_7_31177 = net_31177;
  assign seg_7_14_sp4_r_v_b_9_31179 = net_31179;
  assign seg_7_14_sp4_v_b_6_27746 = net_27746;
  assign seg_7_15_lutff_2_out_27993 = net_27993;
  assign seg_7_15_neigh_op_bnr_6_31399 = seg_8_14_lutff_6_out_31399;
  assign seg_7_15_neigh_op_top_0_28093 = seg_7_16_lutff_0_out_28093;
  assign seg_7_15_sp12_v_b_2_30296 = seg_7_9_sp12_v_b_14_30296;
  assign seg_7_15_sp12_v_b_4_30420 = seg_7_9_sp12_v_b_16_30420;
  assign seg_7_15_sp4_r_v_b_11_31304 = net_31304;
  assign seg_7_15_sp4_r_v_b_31_31546 = net_31546;
  assign seg_7_15_sp4_r_v_b_7_31300 = net_31300;
  assign seg_7_15_sp4_v_b_12_27943 = net_27943;
  assign seg_7_15_sp4_v_b_16_27947 = net_27947;
  assign seg_7_15_sp4_v_b_2_27844 = net_27844;
  assign seg_7_15_sp4_v_b_8_27850 = net_27850;
  assign seg_7_16_lutff_0_out_28093 = net_28093;
  assign seg_7_16_lutff_2_out_28095 = net_28095;
  assign seg_7_16_lutff_3_out_28096 = net_28096;
  assign seg_7_16_lutff_4_out_28097 = net_28097;
  assign seg_7_16_lutff_7_out_28100 = net_28100;
  assign seg_7_16_sp4_v_b_5_27947 = seg_7_15_sp4_v_b_16_27947;
  assign seg_7_17_neigh_op_bot_2_28095 = seg_7_16_lutff_2_out_28095;
  assign seg_7_17_neigh_op_bot_3_28096 = seg_7_16_lutff_3_out_28096;
  assign seg_7_17_neigh_op_bot_4_28097 = seg_7_16_lutff_4_out_28097;
  assign seg_7_17_neigh_op_bot_7_28100 = seg_7_16_lutff_7_out_28100;
  assign seg_7_17_neigh_op_top_0_28297 = seg_7_18_lutff_0_out_28297;
  assign seg_7_17_neigh_op_top_2_28299 = seg_7_18_lutff_2_out_28299;
  assign seg_7_17_neigh_op_top_3_28300 = seg_7_18_lutff_3_out_28300;
  assign seg_7_17_neigh_op_top_5_28302 = seg_7_18_lutff_5_out_28302;
  assign seg_7_17_neigh_op_top_6_28303 = seg_7_18_lutff_6_out_28303;
  assign seg_7_17_sp4_h_l_36_17205 = seg_4_17_sp4_h_r_12_17205;
  assign seg_7_17_sp4_h_r_37_21035 = seg_4_17_sp4_h_r_0_21035;
  assign seg_7_17_sp4_h_r_45_21045 = seg_4_17_sp4_h_r_8_21045;
  assign seg_7_17_sp4_h_r_46_21038 = net_21038;
  assign seg_7_18_lutff_0_out_28297 = net_28297;
  assign seg_7_18_lutff_2_out_28299 = net_28299;
  assign seg_7_18_lutff_3_out_28300 = net_28300;
  assign seg_7_18_lutff_4_out_28301 = net_28301;
  assign seg_7_18_lutff_5_out_28302 = net_28302;
  assign seg_7_18_lutff_6_out_28303 = net_28303;
  assign seg_7_18_neigh_op_top_0_28399 = seg_7_19_lutff_0_out_28399;
  assign seg_7_18_neigh_op_top_3_28402 = seg_7_19_lutff_3_out_28402;
  assign seg_7_18_neigh_op_top_5_28404 = seg_7_19_lutff_5_out_28404;
  assign seg_7_18_neigh_op_top_6_28405 = seg_7_19_lutff_6_out_28405;
  assign seg_7_18_sp4_h_l_37_17327 = seg_5_18_sp4_h_r_24_17327;
  assign seg_7_19_lutff_0_out_28399 = net_28399;
  assign seg_7_19_lutff_3_out_28402 = net_28402;
  assign seg_7_19_lutff_5_out_28404 = net_28404;
  assign seg_7_19_lutff_6_out_28405 = net_28405;
  assign seg_7_19_sp4_h_l_37_17450 = seg_5_19_sp4_h_r_24_17450;
  assign seg_7_1_lutff_1_out_26554 = net_26554;
  assign seg_7_1_sp4_h_l_43_15208 = seg_3_1_sp4_h_r_6_15208;
  assign seg_7_2_lutff_2_out_26631 = net_26631;
  assign seg_7_2_lutff_3_out_26632 = net_26632;
  assign seg_7_2_lutff_4_out_26633 = net_26633;
  assign seg_7_2_sp4_h_l_41_15365 = seg_3_2_sp4_h_r_4_15365;
  assign seg_7_2_sp4_h_l_45_15369 = seg_3_2_sp4_h_r_8_15369;
  assign seg_7_2_sp4_v_b_30_26721 = seg_7_4_sp4_v_b_6_26721;
  assign seg_7_3_lutff_2_out_26769 = net_26769;
  assign seg_7_3_neigh_op_top_0_26869 = seg_7_4_lutff_0_out_26869;
  assign seg_7_3_sp4_h_r_0_30175 = net_30175;
  assign seg_7_3_sp4_h_r_22_26914 = net_26914;
  assign seg_7_3_sp4_h_r_5_30182 = seg_8_3_sp4_h_r_16_30182;
  assign seg_7_3_sp4_h_r_8_30185 = net_30185;
  assign seg_7_4_lutff_0_out_26869 = net_26869;
  assign seg_7_4_lutff_1_out_26870 = net_26870;
  assign seg_7_4_lutff_2_out_26871 = net_26871;
  assign seg_7_4_neigh_op_rgt_4_30167 = seg_8_4_lutff_4_out_30167;
  assign seg_7_4_sp4_h_r_28_23273 = seg_5_4_sp4_h_r_4_23273;
  assign seg_7_4_sp4_h_r_2_30302 = seg_9_4_sp4_h_r_26_30302;
  assign seg_7_4_sp4_h_r_42_19445 = net_19445;
  assign seg_7_4_sp4_h_r_8_30308 = seg_9_4_sp4_h_r_32_30308;
  assign seg_7_4_sp4_r_v_b_27_30189 = net_30189;
  assign seg_7_4_sp4_r_v_b_47_30321 = net_30321;
  assign seg_7_4_sp4_v_b_6_26721 = net_26721;
  assign seg_7_5_lutff_1_out_26972 = net_26972;
  assign seg_7_5_lutff_2_out_26973 = net_26973;
  assign seg_7_5_lutff_3_out_26974 = net_26974;
  assign seg_7_5_lutff_5_out_26976 = net_26976;
  assign seg_7_5_lutff_7_out_26978 = net_26978;
  assign seg_7_5_neigh_op_bot_2_26871 = seg_7_4_lutff_2_out_26871;
  assign seg_7_5_neigh_op_rgt_3_30289 = seg_8_5_lutff_3_out_30289;
  assign seg_7_5_neigh_op_rgt_7_30293 = seg_8_5_lutff_7_out_30293;
  assign seg_7_5_sp4_h_l_36_15729 = seg_4_5_sp4_h_r_12_15729;
  assign seg_7_5_sp4_h_l_42_15737 = seg_4_5_sp4_h_r_18_15737;
  assign seg_7_5_sp4_h_l_44_15739 = seg_4_5_sp4_h_r_20_15739;
  assign seg_7_5_sp4_h_r_10_30423 = seg_9_5_sp4_h_r_34_30423;
  assign seg_7_5_sp4_h_r_22_27118 = seg_9_5_sp4_h_r_46_27118;
  assign seg_7_5_sp4_h_r_24_23390 = net_23390;
  assign seg_7_5_sp4_h_r_47_19561 = seg_4_5_sp4_h_r_10_19561;
  assign seg_7_5_sp4_r_v_b_25_30310 = net_30310;
  assign seg_7_5_sp4_v_b_44_27135 = net_27135;
  assign seg_7_6_lutff_2_out_27075 = net_27075;
  assign seg_7_6_lutff_3_out_27076 = net_27076;
  assign seg_7_6_lutff_7_out_27080 = net_27080;
  assign seg_7_6_neigh_op_bot_1_26972 = seg_7_5_lutff_1_out_26972;
  assign seg_7_6_neigh_op_bot_2_26973 = seg_7_5_lutff_2_out_26973;
  assign seg_7_6_neigh_op_bot_3_26974 = seg_7_5_lutff_3_out_26974;
  assign seg_7_6_neigh_op_bot_5_26976 = seg_7_5_lutff_5_out_26976;
  assign seg_7_6_sp4_h_l_43_15859 = seg_5_6_sp4_h_r_30_15859;
  assign seg_7_6_sp4_h_l_45_15861 = seg_3_6_sp4_h_r_8_15861;
  assign seg_7_6_sp4_h_r_26_23517 = net_23517;
  assign seg_7_6_sp4_h_r_34_23515 = net_23515;
  assign seg_7_6_sp4_h_r_40_19689 = net_19689;
  assign seg_7_6_sp4_h_r_44_19693 = net_19693;
  assign seg_7_6_sp4_v_b_12_27025 = net_27025;
  assign seg_7_6_sp4_v_b_42_27235 = net_27235;
  assign seg_7_7_lutff_0_out_27175 = net_27175;
  assign seg_7_7_lutff_1_out_27176 = net_27176;
  assign seg_7_7_lutff_2_out_27177 = net_27177;
  assign seg_7_7_lutff_3_out_27178 = net_27178;
  assign seg_7_7_lutff_6_out_27181 = net_27181;
  assign seg_7_7_lutff_7_out_27182 = net_27182;
  assign seg_7_7_sp4_h_r_24_23636 = net_23636;
  assign seg_7_7_sp4_h_r_26_23640 = net_23640;
  assign seg_7_7_sp4_v_b_1_27025 = seg_7_6_sp4_v_b_12_27025;
  assign seg_7_7_sp4_v_b_2_27028 = seg_6_4_sp4_r_v_b_39_27028;
  assign seg_7_7_sp4_v_b_6_27032 = seg_6_4_sp4_r_v_b_43_27032;
  assign seg_7_8_lutff_0_out_27277 = net_27277;
  assign seg_7_8_lutff_1_out_27278 = net_27278;
  assign seg_7_8_lutff_2_out_27279 = net_27279;
  assign seg_7_8_lutff_4_out_27281 = net_27281;
  assign seg_7_8_lutff_5_out_27282 = net_27282;
  assign seg_7_8_lutff_6_out_27283 = net_27283;
  assign seg_7_8_lutff_7_out_27284 = net_27284;
  assign seg_7_8_neigh_op_bot_0_27175 = seg_7_7_lutff_0_out_27175;
  assign seg_7_8_neigh_op_bot_6_27181 = seg_7_7_lutff_6_out_27181;
  assign seg_7_8_sp4_h_r_32_23769 = seg_5_8_sp4_h_r_8_23769;
  assign seg_7_8_sp4_h_r_38_19933 = seg_5_8_sp4_h_r_14_19933;
  assign seg_7_8_sp4_h_r_44_19939 = seg_5_8_sp4_h_r_20_19939;
  assign seg_7_8_sp4_v_b_30_27338 = seg_7_10_sp4_v_b_6_27338;
  assign seg_7_8_sp4_v_b_38_27435 = net_27435;
  assign seg_7_8_sp4_v_b_9_27135 = seg_7_5_sp4_v_b_44_27135;
  assign seg_7_9_sp12_v_b_14_30296 = net_30296;
  assign seg_7_9_sp12_v_b_16_30420 = net_30420;
  assign seg_7_9_sp4_h_r_12_27524 = net_27524;
  assign seg_7_9_sp4_h_r_24_23882 = net_23882;
  assign seg_7_9_sp4_r_v_b_38_30927 = seg_8_11_sp4_v_b_14_30927;
  assign seg_7_9_sp4_v_b_34_27444 = net_27444;
  assign seg_7_9_sp4_v_b_36_27535 = net_27535;
  assign seg_7_9_sp4_v_b_38_27537 = net_27537;
  assign seg_7_9_sp4_v_b_7_27235 = seg_7_6_sp4_v_b_42_27235;
  assign seg_8_10_sp4_h_r_4_34873 = seg_10_10_sp4_h_r_28_34873;
  assign seg_8_10_sp4_h_r_8_34877 = seg_10_10_sp4_h_r_32_34877;
  assign seg_8_10_sp4_v_b_34_30936 = net_30936;
  assign seg_8_10_sp4_v_b_36_31048 = net_31048;
  assign seg_8_10_sp4_v_t_37_31172 = seg_7_13_sp4_r_v_b_13_31172;
  assign seg_8_10_sp4_v_t_42_31177 = seg_7_14_sp4_r_v_b_7_31177;
  assign seg_8_11_lutff_0_out_31024 = net_31024;
  assign seg_8_11_lutff_1_out_31025 = net_31025;
  assign seg_8_11_lutff_2_out_31026 = net_31026;
  assign seg_8_11_lutff_3_out_31027 = net_31027;
  assign seg_8_11_lutff_4_out_31028 = net_31028;
  assign seg_8_11_lutff_6_out_31030 = net_31030;
  assign seg_8_11_sp12_v_b_0_33605 = seg_8_5_sp12_v_b_12_33605;
  assign seg_8_11_sp4_h_r_0_34990 = seg_10_11_sp4_h_r_24_34990;
  assign seg_8_11_sp4_h_r_14_31164 = net_31164;
  assign seg_8_11_sp4_h_r_1_34991 = seg_9_11_sp4_h_r_12_34991;
  assign seg_8_11_sp4_h_r_5_34997 = seg_9_11_sp4_h_r_16_34997;
  assign seg_8_11_sp4_h_r_6_34998 = seg_10_11_sp4_h_r_30_34998;
  assign seg_8_11_sp4_r_v_b_15_34759 = net_34759;
  assign seg_8_11_sp4_v_b_10_30813 = net_30813;
  assign seg_8_11_sp4_v_b_14_30927 = net_30927;
  assign seg_8_11_sp4_v_b_26_31051 = seg_8_13_sp4_v_b_2_31051;
  assign seg_8_11_sp4_v_b_44_31179 = seg_7_14_sp4_r_v_b_9_31179;
  assign seg_8_11_sp4_v_t_42_31300 = seg_7_15_sp4_r_v_b_7_31300;
  assign seg_8_11_sp4_v_t_46_31304 = seg_7_15_sp4_r_v_b_11_31304;
  assign seg_8_12_neigh_op_lft_1_27686 = seg_7_12_lutff_1_out_27686;
  assign seg_8_12_neigh_op_lft_2_27687 = seg_7_12_lutff_2_out_27687;
  assign seg_8_12_neigh_op_lft_3_27688 = seg_7_12_lutff_3_out_27688;
  assign seg_8_12_neigh_op_lft_4_27689 = seg_7_12_lutff_4_out_27689;
  assign seg_8_12_neigh_op_lft_5_27690 = seg_7_12_lutff_5_out_27690;
  assign seg_8_12_neigh_op_lft_6_27691 = seg_7_12_lutff_6_out_27691;
  assign seg_8_12_neigh_op_lft_7_27692 = seg_7_12_lutff_7_out_27692;
  assign seg_8_12_neigh_op_rgt_5_34983 = seg_9_12_lutff_5_out_34983;
  assign seg_8_12_neigh_op_tnl_0_27787 = seg_7_13_lutff_0_out_27787;
  assign seg_8_12_sp4_h_l_42_20429 = seg_5_12_sp4_h_r_18_20429;
  assign seg_8_12_sp4_h_l_46_20423 = seg_5_12_sp4_h_r_22_20423;
  assign seg_8_12_sp4_h_r_5_35120 = seg_9_12_sp4_h_r_16_35120;
  assign seg_8_12_sp4_h_r_7_35122 = seg_9_12_sp4_h_r_18_35122;
  assign seg_8_12_sp4_r_v_b_15_34882 = net_34882;
  assign seg_8_12_sp4_v_b_10_30936 = seg_8_10_sp4_v_b_34_30936;
  assign seg_8_13_lutff_0_out_31270 = net_31270;
  assign seg_8_13_lutff_3_out_31273 = net_31273;
  assign seg_8_13_lutff_4_out_31274 = net_31274;
  assign seg_8_13_lutff_5_out_31275 = net_31275;
  assign seg_8_13_lutff_6_out_31276 = net_31276;
  assign seg_8_13_neigh_op_tnl_7_27896 = seg_7_14_lutff_7_out_27896;
  assign seg_8_13_sp4_r_v_b_31_35131 = net_35131;
  assign seg_8_13_sp4_v_b_1_31048 = seg_8_10_sp4_v_b_36_31048;
  assign seg_8_13_sp4_v_b_2_31051 = net_31051;
  assign seg_8_13_sp4_v_b_4_31053 = net_31053;
  assign seg_8_13_sp4_v_t_42_31546 = seg_7_15_sp4_r_v_b_31_31546;
  assign seg_8_14_lutff_0_out_31393 = net_31393;
  assign seg_8_14_lutff_6_out_31399 = net_31399;
  assign seg_8_14_sp4_h_r_7_35368 = seg_11_14_sp4_h_r_42_35368;
  assign seg_8_14_sp4_r_v_b_9_35010 = seg_9_11_sp4_v_b_44_35010;
  assign seg_8_15_neigh_op_bnr_0_35224 = seg_9_14_lutff_0_out_35224;
  assign seg_8_15_neigh_op_rgt_0_35347 = seg_9_15_lutff_0_out_35347;
  assign seg_8_15_neigh_op_rgt_1_35348 = seg_9_15_lutff_1_out_35348;
  assign seg_8_15_neigh_op_rgt_3_35350 = seg_9_15_lutff_3_out_35350;
  assign seg_8_15_neigh_op_rgt_4_35351 = seg_9_15_lutff_4_out_35351;
  assign seg_8_15_neigh_op_rgt_5_35352 = seg_9_15_lutff_5_out_35352;
  assign seg_8_15_neigh_op_rgt_6_35353 = seg_9_15_lutff_6_out_35353;
  assign seg_8_15_neigh_op_rgt_7_35354 = seg_9_15_lutff_7_out_35354;
  assign seg_8_15_sp4_h_r_0_35482 = net_35482;
  assign seg_8_15_sp4_h_r_11_35485 = seg_11_15_sp4_h_r_46_35485;
  assign seg_8_15_sp4_h_r_12_31652 = net_31652;
  assign seg_8_15_sp4_h_r_4_35488 = net_35488;
  assign seg_8_15_sp4_r_v_b_15_35251 = net_35251;
  assign seg_8_15_sp4_r_v_b_39_35497 = net_35497;
  assign seg_8_15_sp4_r_v_b_3_35127 = net_35127;
  assign seg_8_15_sp4_r_v_b_41_35499 = net_35499;
  assign seg_8_15_sp4_r_v_b_4_35130 = seg_9_13_sp4_v_b_28_35130;
  assign seg_8_15_sp4_r_v_b_5_35129 = seg_9_12_sp4_v_b_40_35129;
  assign seg_8_16_sp12_v_b_3_34251 = seg_8_7_sp12_v_b_20_34251;
  assign seg_8_16_sp4_r_v_b_13_35372 = net_35372;
  assign seg_8_16_sp4_r_v_b_19_35378 = net_35378;
  assign seg_8_16_sp4_r_v_b_7_35254 = net_35254;
  assign seg_8_18_sp4_h_l_46_21161 = seg_5_18_sp4_h_r_22_21161;
  assign seg_8_19_sp12_v_t_23_35973 = seg_8_31_span12_vert_0_35973;
  assign seg_8_1_lutff_2_out_29755 = net_29755;
  assign seg_8_1_lutff_3_out_29756 = net_29756;
  assign seg_8_1_lutff_5_out_29758 = net_29758;
  assign seg_8_1_lutff_6_out_29759 = net_29759;
  assign seg_8_1_lutff_7_out_29760 = net_29760;
  assign seg_8_1_neigh_op_lft_1_26554 = seg_7_1_lutff_1_out_26554;
  assign seg_8_1_neigh_op_tnl_2_26631 = seg_7_2_lutff_2_out_26631;
  assign seg_8_1_neigh_op_tnl_4_26633 = seg_7_2_lutff_4_out_26633;
  assign seg_8_21_sp12_v_t_23_36219 = seg_8_31_span12_vert_4_36219;
  assign seg_8_2_lutff_0_out_29881 = net_29881;
  assign seg_8_2_sp4_h_r_4_33889 = net_33889;
  assign seg_8_2_sp4_r_v_b_29_33771 = net_33771;
  assign seg_8_31_span12_vert_0_35973 = net_35973;
  assign seg_8_31_span12_vert_4_36219 = net_36219;
  assign seg_8_3_lutff_5_out_30045 = net_30045;
  assign seg_8_3_lutff_7_out_30047 = net_30047;
  assign seg_8_3_neigh_op_bnr_6_33718 = seg_9_2_lutff_6_out_33718;
  assign seg_8_3_sp4_h_r_16_30182 = net_30182;
  assign seg_8_3_sp4_v_b_28_30069 = net_30069;
  assign seg_8_3_sp4_v_t_36_30310 = seg_7_5_sp4_r_v_b_25_30310;
  assign seg_8_3_sp4_v_t_47_30321 = seg_7_4_sp4_r_v_b_47_30321;
  assign seg_8_4_lutff_2_out_30165 = net_30165;
  assign seg_8_4_lutff_4_out_30167 = net_30167;
  assign seg_8_4_lutff_5_out_30168 = net_30168;
  assign seg_8_4_sp4_h_l_38_19441 = seg_5_4_sp4_h_r_14_19441;
  assign seg_8_4_sp4_h_l_39_19440 = seg_4_4_sp4_h_r_2_19440;
  assign seg_8_4_sp4_h_l_41_19442 = seg_4_4_sp4_h_r_4_19442;
  assign seg_8_4_sp4_h_r_16_30305 = net_30305;
  assign seg_8_4_sp4_h_r_22_30301 = net_30301;
  assign seg_8_4_sp4_r_v_b_13_33896 = net_33896;
  assign seg_8_4_sp4_r_v_b_47_34152 = net_34152;
  assign seg_8_5_lutff_1_out_30287 = net_30287;
  assign seg_8_5_lutff_3_out_30289 = net_30289;
  assign seg_8_5_lutff_4_out_30290 = net_30290;
  assign seg_8_5_lutff_5_out_30291 = net_30291;
  assign seg_8_5_lutff_7_out_30293 = net_30293;
  assign seg_8_5_sp12_v_b_12_33605 = net_33605;
  assign seg_8_5_sp4_h_r_0_34252 = net_34252;
  assign seg_8_5_sp4_h_r_36_23391 = net_23391;
  assign seg_8_5_sp4_h_r_47_23392 = seg_5_5_sp4_h_r_10_23392;
  assign seg_8_5_sp4_v_b_4_30069 = seg_8_3_sp4_v_b_28_30069;
  assign seg_8_6_neigh_op_tnr_1_34364 = seg_9_7_lutff_1_out_34364;
  assign seg_8_6_sp4_r_v_b_19_34148 = net_34148;
  assign seg_8_6_sp4_v_b_22_30320 = net_30320;
  assign seg_8_6_sp4_v_b_26_30436 = net_30436;
  assign seg_8_6_sp4_v_b_30_30440 = net_30440;
  assign seg_8_6_sp4_v_b_32_30442 = net_30442;
  assign seg_8_6_sp4_v_b_3_30189 = seg_7_4_sp4_r_v_b_27_30189;
  assign seg_8_6_sp4_v_b_40_30560 = net_30560;
  assign seg_8_6_sp4_v_b_44_30564 = net_30564;
  assign seg_8_7_sp12_v_b_20_34251 = net_34251;
  assign seg_8_7_sp4_h_l_41_19811 = seg_4_7_sp4_h_r_4_19811;
  assign seg_8_7_sp4_h_l_42_19814 = seg_5_7_sp4_h_r_18_19814;
  assign seg_8_7_sp4_h_r_0_34498 = seg_10_7_sp4_h_r_24_34498;
  assign seg_8_7_sp4_h_r_7_34507 = seg_9_7_sp4_h_r_18_34507;
  assign seg_8_7_sp4_r_v_b_29_34391 = net_34391;
  assign seg_8_7_sp4_v_b_11_30320 = seg_8_6_sp4_v_b_22_30320;
  assign seg_8_7_sp4_v_b_32_30565 = net_30565;
  assign seg_8_8_lutff_1_out_30656 = net_30656;
  assign seg_8_8_lutff_2_out_30657 = net_30657;
  assign seg_8_8_lutff_3_out_30658 = net_30658;
  assign seg_8_8_lutff_4_out_30659 = net_30659;
  assign seg_8_8_lutff_5_out_30660 = net_30660;
  assign seg_8_8_lutff_6_out_30661 = net_30661;
  assign seg_8_8_lutff_7_out_30662 = net_30662;
  assign seg_8_8_neigh_op_bnl_1_27176 = seg_7_7_lutff_1_out_27176;
  assign seg_8_8_neigh_op_lft_1_27278 = seg_7_8_lutff_1_out_27278;
  assign seg_8_8_neigh_op_lft_2_27279 = seg_7_8_lutff_2_out_27279;
  assign seg_8_8_neigh_op_lft_4_27281 = seg_7_8_lutff_4_out_27281;
  assign seg_8_8_neigh_op_lft_5_27282 = seg_7_8_lutff_5_out_27282;
  assign seg_8_8_neigh_op_lft_6_27283 = seg_7_8_lutff_6_out_27283;
  assign seg_8_8_neigh_op_lft_7_27284 = seg_7_8_lutff_7_out_27284;
  assign seg_8_8_neigh_op_tnr_1_34610 = seg_9_9_lutff_1_out_34610;
  assign seg_8_8_neigh_op_tnr_2_34611 = seg_9_9_lutff_2_out_34611;
  assign seg_8_8_neigh_op_tnr_4_34613 = seg_9_9_lutff_4_out_34613;
  assign seg_8_8_neigh_op_top_4_30782 = seg_8_9_lutff_4_out_30782;
  assign seg_8_8_neigh_op_top_5_30783 = seg_8_9_lutff_5_out_30783;
  assign seg_8_8_neigh_op_top_7_30785 = seg_8_9_lutff_7_out_30785;
  assign seg_8_8_sp4_h_r_11_34624 = seg_11_8_sp4_h_r_46_34624;
  assign seg_8_8_sp4_h_r_3_34626 = seg_11_8_sp4_h_r_38_34626;
  assign seg_8_8_sp4_h_r_7_34630 = seg_11_8_sp4_h_r_42_34630;
  assign seg_8_8_sp4_h_r_9_34632 = seg_11_8_sp4_h_r_44_34632;
  assign seg_8_8_sp4_v_b_2_30436 = seg_8_6_sp4_v_b_26_30436;
  assign seg_8_8_sp4_v_b_47_30813 = seg_8_11_sp4_v_b_10_30813;
  assign seg_8_8_sp4_v_b_6_30440 = seg_8_6_sp4_v_b_30_30440;
  assign seg_8_8_sp4_v_b_8_30442 = seg_8_6_sp4_v_b_32_30442;
  assign seg_8_9_lutff_1_out_30779 = net_30779;
  assign seg_8_9_lutff_2_out_30780 = net_30780;
  assign seg_8_9_lutff_4_out_30782 = net_30782;
  assign seg_8_9_lutff_5_out_30783 = net_30783;
  assign seg_8_9_lutff_6_out_30784 = net_30784;
  assign seg_8_9_lutff_7_out_30785 = net_30785;
  assign seg_8_9_neigh_op_tnl_2_27483 = seg_7_10_lutff_2_out_27483;
  assign seg_8_9_neigh_op_tnl_4_27485 = seg_7_10_lutff_4_out_27485;
  assign seg_8_9_sp4_r_v_b_1_34387 = net_34387;
  assign seg_8_9_sp4_v_b_5_30560 = seg_8_6_sp4_v_b_40_30560;
  assign seg_8_9_sp4_v_b_8_30565 = seg_8_7_sp4_v_b_32_30565;
  assign seg_8_9_sp4_v_b_9_30564 = seg_8_6_sp4_v_b_44_30564;
  assign seg_8_9_sp4_v_t_41_31053 = seg_8_13_sp4_v_b_4_31053;
  assign seg_9_10_lutff_1_out_34733 = net_34733;
  assign seg_9_10_lutff_2_out_34734 = net_34734;
  assign seg_9_10_lutff_4_out_34736 = net_34736;
  assign seg_9_10_lutff_5_out_34737 = net_34737;
  assign seg_9_10_lutff_6_out_34738 = net_34738;
  assign seg_9_10_neigh_op_tnl_4_31028 = seg_8_11_lutff_4_out_31028;
  assign seg_9_10_sp4_h_r_11_38701 = seg_12_10_sp4_h_r_46_38701;
  assign seg_9_10_sp4_h_r_3_38703 = seg_10_10_sp4_h_r_14_38703;
  assign seg_9_10_sp4_r_v_b_31_38593 = net_38593;
  assign seg_9_10_sp4_v_b_0_34511 = net_34511;
  assign seg_9_10_sp4_v_b_46_34889 = net_34889;
  assign seg_9_11_lutff_0_out_34855 = net_34855;
  assign seg_9_11_lutff_6_out_34861 = net_34861;
  assign seg_9_11_sp4_h_r_12_34991 = net_34991;
  assign seg_9_11_sp4_h_r_16_34997 = net_34997;
  assign seg_9_11_sp4_h_r_28_31165 = net_31165;
  assign seg_9_11_sp4_h_r_32_31169 = net_31169;
  assign seg_9_11_sp4_h_r_44_27738 = net_27738;
  assign seg_9_11_sp4_r_v_b_13_38588 = net_38588;
  assign seg_9_11_sp4_r_v_b_17_38592 = net_38592;
  assign seg_9_11_sp4_r_v_b_1_38464 = net_38464;
  assign seg_9_11_sp4_v_b_0_34634 = net_34634;
  assign seg_9_11_sp4_v_b_12_34756 = net_34756;
  assign seg_9_11_sp4_v_b_16_34760 = net_34760;
  assign seg_9_11_sp4_v_b_28_34884 = net_34884;
  assign seg_9_11_sp4_v_b_44_35010 = net_35010;
  assign seg_9_11_sp4_v_t_38_35127 = seg_8_15_sp4_r_v_b_3_35127;
  assign seg_9_11_sp4_v_t_42_35131 = seg_8_13_sp4_r_v_b_31_35131;
  assign seg_9_12_lutff_5_out_34983 = net_34983;
  assign seg_9_12_neigh_op_bnl_3_31027 = seg_8_11_lutff_3_out_31027;
  assign seg_9_12_neigh_op_tnl_5_31275 = seg_8_13_lutff_5_out_31275;
  assign seg_9_12_sp12_v_b_1_37438 = seg_9_7_sp12_v_b_10_37438;
  assign seg_9_12_sp4_h_r_16_35120 = net_35120;
  assign seg_9_12_sp4_h_r_18_35122 = net_35122;
  assign seg_9_12_sp4_h_r_9_38955 = seg_10_12_sp4_h_r_20_38955;
  assign seg_9_12_sp4_r_v_b_22_38720 = seg_10_10_sp4_v_b_46_38720;
  assign seg_9_12_sp4_v_b_1_34756 = seg_9_11_sp4_v_b_12_34756;
  assign seg_9_12_sp4_v_b_40_35129 = net_35129;
  assign seg_9_12_sp4_v_t_39_35251 = seg_8_15_sp4_r_v_b_15_35251;
  assign seg_9_12_sp4_v_t_42_35254 = seg_8_16_sp4_r_v_b_7_35254;
  assign seg_9_13_lutff_3_out_35104 = net_35104;
  assign seg_9_13_neigh_op_rgt_1_38933 = seg_10_13_lutff_1_out_38933;
  assign seg_9_13_sp12_h_r_3_35232 = seg_14_13_sp12_h_r_12_35232;
  assign seg_9_13_sp4_h_r_10_39069 = net_39069;
  assign seg_9_13_sp4_h_r_1_39068 = seg_12_13_sp4_h_r_36_39068;
  assign seg_9_13_sp4_v_b_11_34889 = seg_9_10_sp4_v_b_46_34889;
  assign seg_9_13_sp4_v_b_28_35130 = net_35130;
  assign seg_9_13_sp4_v_b_4_34884 = seg_9_11_sp4_v_b_28_34884;
  assign seg_9_13_sp4_v_t_37_35372 = seg_8_16_sp4_r_v_b_13_35372;
  assign seg_9_13_sp4_v_t_43_35378 = seg_8_16_sp4_r_v_b_19_35378;
  assign seg_9_14_lutff_0_out_35224 = net_35224;
  assign seg_9_14_lutff_2_out_35226 = net_35226;
  assign seg_9_14_lutff_3_out_35227 = net_35227;
  assign seg_9_14_lutff_4_out_35228 = net_35228;
  assign seg_9_14_lutff_7_out_35231 = net_35231;
  assign seg_9_14_neigh_op_bnr_2_38934 = seg_10_13_lutff_2_out_38934;
  assign seg_9_14_sp4_h_r_26_31532 = net_31532;
  assign seg_9_14_sp4_h_r_5_39197 = seg_10_14_sp4_h_r_16_39197;
  assign seg_9_14_sp4_v_b_9_35010 = seg_9_11_sp4_v_b_44_35010;
  assign seg_9_14_sp4_v_t_39_35497 = seg_8_15_sp4_r_v_b_39_35497;
  assign seg_9_14_sp4_v_t_41_35499 = seg_8_15_sp4_r_v_b_41_35499;
  assign seg_9_15_lutff_0_out_35347 = net_35347;
  assign seg_9_15_lutff_1_out_35348 = net_35348;
  assign seg_9_15_lutff_3_out_35350 = net_35350;
  assign seg_9_15_lutff_4_out_35351 = net_35351;
  assign seg_9_15_lutff_5_out_35352 = net_35352;
  assign seg_9_15_lutff_6_out_35353 = net_35353;
  assign seg_9_15_lutff_7_out_35354 = net_35354;
  assign seg_9_15_neigh_op_bot_4_35228 = seg_9_14_lutff_4_out_35228;
  assign seg_9_15_neigh_op_bot_7_35231 = seg_9_14_lutff_7_out_35231;
  assign seg_9_15_neigh_op_rgt_0_39178 = seg_10_15_lutff_0_out_39178;
  assign seg_9_15_neigh_op_rgt_4_39182 = seg_10_15_lutff_4_out_39182;
  assign seg_9_15_sp4_h_r_36_28136 = net_28136;
  assign seg_9_15_sp4_h_r_3_39318 = seg_12_15_sp4_h_r_38_39318;
  assign seg_9_16_sp4_h_r_0_39436 = net_39436;
  assign seg_9_16_sp4_r_v_b_31_39331 = net_39331;
  assign seg_9_16_sp4_r_v_b_41_39453 = net_39453;
  assign seg_9_16_sp4_r_v_b_43_39455 = net_39455;
  assign seg_9_16_sp4_v_b_38_35619 = net_35619;
  assign seg_9_17_lutff_0_out_35593 = net_35593;
  assign seg_9_17_lutff_2_out_35595 = net_35595;
  assign seg_9_17_lutff_3_out_35596 = net_35596;
  assign seg_9_17_neigh_op_bnr_1_39302 = seg_10_16_lutff_1_out_39302;
  assign seg_9_17_neigh_op_bnr_3_39304 = seg_10_16_lutff_3_out_39304;
  assign seg_9_17_sp4_h_l_39_24870 = seg_5_17_sp4_h_r_2_24870;
  assign seg_9_17_sp4_r_v_b_35_39458 = net_39458;
  assign seg_9_18_lutff_0_out_35716 = net_35716;
  assign seg_9_18_lutff_2_out_35718 = net_35718;
  assign seg_9_18_lutff_5_out_35721 = net_35721;
  assign seg_9_18_lutff_6_out_35722 = net_35722;
  assign seg_9_18_lutff_7_out_35723 = net_35723;
  assign seg_9_18_neigh_op_bnr_0_39424 = seg_10_17_lutff_0_out_39424;
  assign seg_9_18_neigh_op_bnr_1_39425 = seg_10_17_lutff_1_out_39425;
  assign seg_9_18_neigh_op_bnr_2_39426 = seg_10_17_lutff_2_out_39426;
  assign seg_9_18_neigh_op_bnr_4_39428 = seg_10_17_lutff_4_out_39428;
  assign seg_9_18_neigh_op_bnr_6_39430 = seg_10_17_lutff_6_out_39430;
  assign seg_9_18_neigh_op_bnr_7_39431 = seg_10_17_lutff_7_out_39431;
  assign seg_9_18_neigh_op_bot_2_35595 = seg_9_17_lutff_2_out_35595;
  assign seg_9_18_sp4_r_v_b_17_39453 = seg_9_16_sp4_r_v_b_41_39453;
  assign seg_9_18_sp4_r_v_b_19_39455 = seg_9_16_sp4_r_v_b_43_39455;
  assign seg_9_18_sp4_r_v_b_1_39325 = seg_10_15_sp4_v_b_36_39325;
  assign seg_9_18_sp4_r_v_b_22_39458 = seg_9_17_sp4_r_v_b_35_39458;
  assign seg_9_18_sp4_r_v_b_35_39581 = net_39581;
  assign seg_9_18_sp4_r_v_b_7_39331 = seg_9_16_sp4_r_v_b_31_39331;
  assign seg_9_18_sp4_v_b_14_35619 = seg_9_16_sp4_v_b_38_35619;
  assign seg_9_1_lutff_1_out_33585 = net_33585;
  assign seg_9_1_lutff_3_out_33587 = net_33587;
  assign seg_9_1_lutff_4_out_33588 = net_33588;
  assign seg_9_1_lutff_6_out_33590 = net_33590;
  assign seg_9_1_lutff_7_out_33591 = net_33591;
  assign seg_9_1_neigh_op_lft_3_29756 = seg_8_1_lutff_3_out_29756;
  assign seg_9_1_neigh_op_lft_5_29758 = seg_8_1_lutff_5_out_29758;
  assign seg_9_1_neigh_op_lft_7_29760 = seg_8_1_lutff_7_out_29760;
  assign seg_9_1_sp4_v_t_37_33896 = seg_8_4_sp4_r_v_b_13_33896;
  assign seg_9_1_sp4_v_t_45_33904 = seg_9_5_sp4_v_b_8_33904;
  assign seg_9_2_lutff_3_out_33715 = net_33715;
  assign seg_9_2_lutff_6_out_33718 = net_33718;
  assign seg_9_2_sp4_h_r_3_37719 = seg_12_2_sp4_h_r_38_37719;
  assign seg_9_3_lutff_3_out_33874 = net_33874;
  assign seg_9_3_neigh_op_bot_3_33715 = seg_9_2_lutff_3_out_33715;
  assign seg_9_3_sp4_h_r_5_37844 = seg_12_3_sp4_h_r_40_37844;
  assign seg_9_3_sp4_v_b_28_33900 = net_33900;
  assign seg_9_3_sp4_v_t_47_34152 = seg_8_4_sp4_r_v_b_47_34152;
  assign seg_9_4_lutff_2_out_33996 = net_33996;
  assign seg_9_4_lutff_6_out_34000 = net_34000;
  assign seg_9_4_lutff_7_out_34001 = net_34001;
  assign seg_9_4_neigh_op_rgt_3_37828 = seg_10_4_lutff_3_out_37828;
  assign seg_9_4_sp4_h_r_26_30302 = net_30302;
  assign seg_9_4_sp4_h_r_32_30308 = net_30308;
  assign seg_9_4_sp4_v_b_5_33771 = seg_8_2_sp4_r_v_b_29_33771;
  assign seg_9_5_lutff_0_out_34117 = net_34117;
  assign seg_9_5_lutff_3_out_34120 = net_34120;
  assign seg_9_5_lutff_6_out_34123 = net_34123;
  assign seg_9_5_sp4_h_r_34_30423 = net_30423;
  assign seg_9_5_sp4_h_r_46_27118 = net_27118;
  assign seg_9_5_sp4_v_b_4_33900 = seg_9_3_sp4_v_b_28_33900;
  assign seg_9_5_sp4_v_b_8_33904 = net_33904;
  assign seg_9_5_sp4_v_t_36_34387 = seg_8_9_sp4_r_v_b_1_34387;
  assign seg_9_5_sp4_v_t_38_34389 = seg_9_8_sp4_v_b_14_34389;
  assign seg_9_6_lutff_0_out_34240 = net_34240;
  assign seg_9_6_lutff_2_out_34242 = net_34242;
  assign seg_9_6_neigh_op_top_7_34370 = seg_9_7_lutff_7_out_34370;
  assign seg_9_6_sp4_h_r_22_34378 = net_34378;
  assign seg_9_6_sp4_h_r_5_38213 = seg_12_6_sp4_h_r_40_38213;
  assign seg_9_6_sp4_r_v_b_9_37857 = net_37857;
  assign seg_9_6_sp4_v_t_36_34510 = seg_9_9_sp4_v_b_12_34510;
  assign seg_9_7_lutff_0_out_34363 = net_34363;
  assign seg_9_7_lutff_1_out_34364 = net_34364;
  assign seg_9_7_lutff_2_out_34365 = net_34365;
  assign seg_9_7_lutff_3_out_34366 = net_34366;
  assign seg_9_7_lutff_4_out_34367 = net_34367;
  assign seg_9_7_lutff_6_out_34369 = net_34369;
  assign seg_9_7_lutff_7_out_34370 = net_34370;
  assign seg_9_7_neigh_op_top_1_34487 = seg_9_8_lutff_1_out_34487;
  assign seg_9_7_sp12_h_r_18_1555 = net_1555;
  assign seg_9_7_sp12_h_r_1_38326 = seg_18_7_sp12_h_r_18_38326;
  assign seg_9_7_sp12_v_b_10_37438 = net_37438;
  assign seg_9_7_sp4_h_r_18_34507 = net_34507;
  assign seg_9_7_sp4_r_v_b_35_38228 = net_38228;
  assign seg_9_7_sp4_r_v_b_3_37974 = net_37974;
  assign seg_9_7_sp4_v_b_37_34511 = seg_9_10_sp4_v_b_0_34511;
  assign seg_9_7_sp4_v_b_6_34148 = seg_8_6_sp4_r_v_b_19_34148;
  assign seg_9_7_sp4_v_t_37_34634 = seg_9_11_sp4_v_b_0_34634;
  assign seg_9_7_sp4_v_t_43_34640 = seg_9_9_sp4_v_b_30_34640;
  assign seg_9_8_lutff_1_out_34487 = net_34487;
  assign seg_9_8_lutff_2_out_34488 = net_34488;
  assign seg_9_8_lutff_3_out_34489 = net_34489;
  assign seg_9_8_lutff_4_out_34490 = net_34490;
  assign seg_9_8_lutff_5_out_34491 = net_34491;
  assign seg_9_8_lutff_6_out_34492 = net_34492;
  assign seg_9_8_neigh_op_lft_1_30656 = seg_8_8_lutff_1_out_30656;
  assign seg_9_8_neigh_op_lft_2_30657 = seg_8_8_lutff_2_out_30657;
  assign seg_9_8_neigh_op_lft_3_30658 = seg_8_8_lutff_3_out_30658;
  assign seg_9_8_neigh_op_lft_4_30659 = seg_8_8_lutff_4_out_30659;
  assign seg_9_8_neigh_op_lft_5_30660 = seg_8_8_lutff_5_out_30660;
  assign seg_9_8_neigh_op_lft_6_30661 = seg_8_8_lutff_6_out_30661;
  assign seg_9_8_neigh_op_lft_7_30662 = seg_8_8_lutff_7_out_30662;
  assign seg_9_8_neigh_op_tnl_1_30779 = seg_8_9_lutff_1_out_30779;
  assign seg_9_8_sp4_h_l_43_23767 = seg_5_8_sp4_h_r_6_23767;
  assign seg_9_8_sp4_h_r_30_30798 = net_30798;
  assign seg_9_8_sp4_v_b_14_34389 = net_34389;
  assign seg_9_8_sp4_v_t_36_34756 = seg_9_11_sp4_v_b_12_34756;
  assign seg_9_8_sp4_v_t_39_34759 = seg_8_11_sp4_r_v_b_15_34759;
  assign seg_9_8_sp4_v_t_40_34760 = seg_9_11_sp4_v_b_16_34760;
  assign seg_9_9_lutff_0_out_34609 = net_34609;
  assign seg_9_9_lutff_1_out_34610 = net_34610;
  assign seg_9_9_lutff_2_out_34611 = net_34611;
  assign seg_9_9_lutff_3_out_34612 = net_34612;
  assign seg_9_9_lutff_4_out_34613 = net_34613;
  assign seg_9_9_lutff_5_out_34614 = net_34614;
  assign seg_9_9_neigh_op_top_2_34734 = seg_9_10_lutff_2_out_34734;
  assign seg_9_9_neigh_op_top_5_34737 = seg_9_10_lutff_5_out_34737;
  assign seg_9_9_neigh_op_top_6_34738 = seg_9_10_lutff_6_out_34738;
  assign seg_9_9_sp4_v_b_12_34510 = net_34510;
  assign seg_9_9_sp4_v_b_30_34640 = net_34640;
  assign seg_9_9_sp4_v_b_5_34391 = seg_8_7_sp4_r_v_b_29_34391;
  assign seg_9_9_sp4_v_t_39_34882 = seg_8_12_sp4_r_v_b_15_34882;
  wire gnd, vcc;
  GND gnd_cell (.Y(gnd));
  VCC vcc_cell (.Y(vcc));
  inout io_4_31_0;
  wire io_pad_4_31_0_din;
  wire io_pad_4_31_0_dout;
  wire io_pad_4_31_0_oe;
  IO_PAD io_pad_4_31_0 (
    .DIN(io_pad_4_31_0_din),
    .DOUT(io_pad_4_31_0_dout),
    .OE(io_pad_4_31_0_oe),
    .PACKAGEPIN(io_4_31_0)
  );
  inout io_5_31_0;
  wire io_pad_5_31_0_din;
  wire io_pad_5_31_0_dout;
  wire io_pad_5_31_0_oe;
  IO_PAD io_pad_5_31_0 (
    .DIN(io_pad_5_31_0_din),
    .DOUT(io_pad_5_31_0_dout),
    .OE(io_pad_5_31_0_oe),
    .PACKAGEPIN(io_5_31_0)
  );
  inout io_5_0_0;
  wire io_pad_5_0_0_din;
  wire io_pad_5_0_0_dout;
  wire io_pad_5_0_0_oe;
  IO_PAD io_pad_5_0_0 (
    .DIN(io_pad_5_0_0_din),
    .DOUT(io_pad_5_0_0_dout),
    .OE(io_pad_5_0_0_oe),
    .PACKAGEPIN(io_5_0_0)
  );
  inout io_6_0_0;
  wire io_pad_6_0_0_din;
  wire io_pad_6_0_0_dout;
  wire io_pad_6_0_0_oe;
  IO_PAD io_pad_6_0_0 (
    .DIN(io_pad_6_0_0_din),
    .DOUT(io_pad_6_0_0_dout),
    .OE(io_pad_6_0_0_oe),
    .PACKAGEPIN(io_6_0_0)
  );
  inout io_6_0_1;
  wire io_pad_6_0_1_din;
  wire io_pad_6_0_1_dout;
  wire io_pad_6_0_1_oe;
  IO_PAD io_pad_6_0_1 (
    .DIN(io_pad_6_0_1_din),
    .DOUT(io_pad_6_0_1_dout),
    .OE(io_pad_6_0_1_oe),
    .PACKAGEPIN(io_6_0_1)
  );
  inout io_6_31_0;
  wire io_pad_6_31_0_din;
  wire io_pad_6_31_0_dout;
  wire io_pad_6_31_0_oe;
  IO_PAD io_pad_6_31_0 (
    .DIN(io_pad_6_31_0_din),
    .DOUT(io_pad_6_31_0_dout),
    .OE(io_pad_6_31_0_oe),
    .PACKAGEPIN(io_6_31_0)
  );
  inout io_7_0_0;
  wire io_pad_7_0_0_din;
  wire io_pad_7_0_0_dout;
  wire io_pad_7_0_0_oe;
  IO_PAD io_pad_7_0_0 (
    .DIN(io_pad_7_0_0_din),
    .DOUT(io_pad_7_0_0_dout),
    .OE(io_pad_7_0_0_oe),
    .PACKAGEPIN(io_7_0_0)
  );
  inout io_8_31_0;
  wire io_pad_8_31_0_din;
  wire io_pad_8_31_0_dout;
  wire io_pad_8_31_0_oe;
  IO_PAD io_pad_8_31_0 (
    .DIN(io_pad_8_31_0_din),
    .DOUT(io_pad_8_31_0_dout),
    .OE(io_pad_8_31_0_oe),
    .PACKAGEPIN(io_8_31_0)
  );
  inout io_8_31_1;
  wire io_pad_8_31_1_din;
  wire io_pad_8_31_1_dout;
  wire io_pad_8_31_1_oe;
  IO_PAD io_pad_8_31_1 (
    .DIN(io_pad_8_31_1_din),
    .DOUT(io_pad_8_31_1_dout),
    .OE(io_pad_8_31_1_oe),
    .PACKAGEPIN(io_8_31_1)
  );
  inout io_8_0_0;
  wire io_pad_8_0_0_din;
  wire io_pad_8_0_0_dout;
  wire io_pad_8_0_0_oe;
  IO_PAD io_pad_8_0_0 (
    .DIN(io_pad_8_0_0_din),
    .DOUT(io_pad_8_0_0_dout),
    .OE(io_pad_8_0_0_oe),
    .PACKAGEPIN(io_8_0_0)
  );
  inout io_9_0_0;
  wire io_pad_9_0_0_din;
  wire io_pad_9_0_0_dout;
  wire io_pad_9_0_0_oe;
  IO_PAD io_pad_9_0_0 (
    .DIN(io_pad_9_0_0_din),
    .DOUT(io_pad_9_0_0_dout),
    .OE(io_pad_9_0_0_oe),
    .PACKAGEPIN(io_9_0_0)
  );
  inout io_9_0_1;
  wire io_pad_9_0_1_din;
  wire io_pad_9_0_1_dout;
  wire io_pad_9_0_1_oe;
  IO_PAD io_pad_9_0_1 (
    .DIN(io_pad_9_0_1_din),
    .DOUT(io_pad_9_0_1_dout),
    .OE(io_pad_9_0_1_oe),
    .PACKAGEPIN(io_9_0_1)
  );
  inout io_12_31_1;
  wire io_pad_12_31_1_din;
  wire io_pad_12_31_1_dout;
  wire io_pad_12_31_1_oe;
  IO_PAD io_pad_12_31_1 (
    .DIN(io_pad_12_31_1_din),
    .DOUT(io_pad_12_31_1_dout),
    .OE(io_pad_12_31_1_oe),
    .PACKAGEPIN(io_12_31_1)
  );
  inout io_13_0_1;
  wire io_pad_13_0_1_din;
  wire io_pad_13_0_1_dout;
  wire io_pad_13_0_1_oe;
  IO_PAD io_pad_13_0_1 (
    .DIN(io_pad_13_0_1_din),
    .DOUT(io_pad_13_0_1_dout),
    .OE(io_pad_13_0_1_oe),
    .PACKAGEPIN(io_13_0_1)
  );
  inout io_13_31_0;
  wire io_pad_13_31_0_din;
  wire io_pad_13_31_0_dout;
  wire io_pad_13_31_0_oe;
  IO_PAD io_pad_13_31_0 (
    .DIN(io_pad_13_31_0_din),
    .DOUT(io_pad_13_31_0_dout),
    .OE(io_pad_13_31_0_oe),
    .PACKAGEPIN(io_13_31_0)
  );
  inout io_13_31_1;
  wire io_pad_13_31_1_din;
  wire io_pad_13_31_1_dout;
  wire io_pad_13_31_1_oe;
  IO_PAD io_pad_13_31_1 (
    .DIN(io_pad_13_31_1_din),
    .DOUT(io_pad_13_31_1_dout),
    .OE(io_pad_13_31_1_oe),
    .PACKAGEPIN(io_13_31_1)
  );
  inout io_15_0_0;
  wire io_pad_15_0_0_din;
  wire io_pad_15_0_0_dout;
  wire io_pad_15_0_0_oe;
  IO_PAD io_pad_15_0_0 (
    .DIN(io_pad_15_0_0_din),
    .DOUT(io_pad_15_0_0_dout),
    .OE(io_pad_15_0_0_oe),
    .PACKAGEPIN(io_15_0_0)
  );
  inout io_16_0_0;
  wire io_pad_16_0_0_din;
  wire io_pad_16_0_0_dout;
  wire io_pad_16_0_0_oe;
  IO_PAD io_pad_16_0_0 (
    .DIN(io_pad_16_0_0_din),
    .DOUT(io_pad_16_0_0_dout),
    .OE(io_pad_16_0_0_oe),
    .PACKAGEPIN(io_16_0_0)
  );
  inout io_17_0_0;
  wire io_pad_17_0_0_din;
  wire io_pad_17_0_0_dout;
  wire io_pad_17_0_0_oe;
  IO_PAD io_pad_17_0_0 (
    .DIN(io_pad_17_0_0_din),
    .DOUT(io_pad_17_0_0_dout),
    .OE(io_pad_17_0_0_oe),
    .PACKAGEPIN(io_17_0_0)
  );
  inout io_16_31_0;
  wire io_pad_16_31_0_din;
  wire io_pad_16_31_0_dout;
  wire io_pad_16_31_0_oe;
  IO_PAD io_pad_16_31_0 (
    .DIN(io_pad_16_31_0_din),
    .DOUT(io_pad_16_31_0_dout),
    .OE(io_pad_16_31_0_oe),
    .PACKAGEPIN(io_16_31_0)
  );
  inout io_16_31_1;
  wire io_pad_16_31_1_din;
  wire io_pad_16_31_1_dout;
  wire io_pad_16_31_1_oe;
  IO_PAD io_pad_16_31_1 (
    .DIN(io_pad_16_31_1_din),
    .DOUT(io_pad_16_31_1_dout),
    .OE(io_pad_16_31_1_oe),
    .PACKAGEPIN(io_16_31_1)
  );
  inout io_18_0_0;
  wire io_pad_18_0_0_din;
  wire io_pad_18_0_0_dout;
  wire io_pad_18_0_0_oe;
  IO_PAD io_pad_18_0_0 (
    .DIN(io_pad_18_0_0_din),
    .DOUT(io_pad_18_0_0_dout),
    .OE(io_pad_18_0_0_oe),
    .PACKAGEPIN(io_18_0_0)
  );
  inout io_17_31_0;
  wire io_pad_17_31_0_din;
  wire io_pad_17_31_0_dout;
  wire io_pad_17_31_0_oe;
  IO_PAD io_pad_17_31_0 (
    .DIN(io_pad_17_31_0_din),
    .DOUT(io_pad_17_31_0_dout),
    .OE(io_pad_17_31_0_oe),
    .PACKAGEPIN(io_17_31_0)
  );
  inout io_18_0_1;
  wire io_pad_18_0_1_din;
  wire io_pad_18_0_1_dout;
  wire io_pad_18_0_1_oe;
  IO_PAD io_pad_18_0_1 (
    .DIN(io_pad_18_0_1_din),
    .DOUT(io_pad_18_0_1_dout),
    .OE(io_pad_18_0_1_oe),
    .PACKAGEPIN(io_18_0_1)
  );
  inout io_19_0_0;
  wire io_pad_19_0_0_din;
  wire io_pad_19_0_0_dout;
  wire io_pad_19_0_0_oe;
  IO_PAD io_pad_19_0_0 (
    .DIN(io_pad_19_0_0_din),
    .DOUT(io_pad_19_0_0_dout),
    .OE(io_pad_19_0_0_oe),
    .PACKAGEPIN(io_19_0_0)
  );
  inout io_19_0_1;
  wire io_pad_19_0_1_din;
  wire io_pad_19_0_1_dout;
  wire io_pad_19_0_1_oe;
  IO_PAD io_pad_19_0_1 (
    .DIN(io_pad_19_0_1_din),
    .DOUT(io_pad_19_0_1_dout),
    .OE(io_pad_19_0_1_oe),
    .PACKAGEPIN(io_19_0_1)
  );
  inout io_18_31_0;
  wire io_pad_18_31_0_din;
  wire io_pad_18_31_0_dout;
  wire io_pad_18_31_0_oe;
  IO_PAD io_pad_18_31_0 (
    .DIN(io_pad_18_31_0_din),
    .DOUT(io_pad_18_31_0_dout),
    .OE(io_pad_18_31_0_oe),
    .PACKAGEPIN(io_18_31_0)
  );
  inout io_18_31_1;
  wire io_pad_18_31_1_din;
  wire io_pad_18_31_1_dout;
  wire io_pad_18_31_1_oe;
  IO_PAD io_pad_18_31_1 (
    .DIN(io_pad_18_31_1_din),
    .DOUT(io_pad_18_31_1_dout),
    .OE(io_pad_18_31_1_oe),
    .PACKAGEPIN(io_18_31_1)
  );
  inout io_21_0_1;
  wire io_pad_21_0_1_din;
  wire io_pad_21_0_1_dout;
  wire io_pad_21_0_1_oe;
  IO_PAD io_pad_21_0_1 (
    .DIN(io_pad_21_0_1_din),
    .DOUT(io_pad_21_0_1_dout),
    .OE(io_pad_21_0_1_oe),
    .PACKAGEPIN(io_21_0_1)
  );
  inout io_22_0_1;
  wire io_pad_22_0_1_din;
  wire io_pad_22_0_1_dout;
  wire io_pad_22_0_1_oe;
  IO_PAD io_pad_22_0_1 (
    .DIN(io_pad_22_0_1_din),
    .DOUT(io_pad_22_0_1_dout),
    .OE(io_pad_22_0_1_oe),
    .PACKAGEPIN(io_22_0_1)
  );
  inout io_23_0_0;
  wire io_pad_23_0_0_din;
  wire io_pad_23_0_0_dout;
  wire io_pad_23_0_0_oe;
  IO_PAD io_pad_23_0_0 (
    .DIN(io_pad_23_0_0_din),
    .DOUT(io_pad_23_0_0_dout),
    .OE(io_pad_23_0_0_oe),
    .PACKAGEPIN(io_23_0_0)
  );
  inout io_23_0_1;
  wire io_pad_23_0_1_din;
  wire io_pad_23_0_1_dout;
  wire io_pad_23_0_1_oe;
  IO_PAD io_pad_23_0_1 (
    .DIN(io_pad_23_0_1_din),
    .DOUT(io_pad_23_0_1_dout),
    .OE(io_pad_23_0_1_oe),
    .PACKAGEPIN(io_23_0_1)
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_0_10_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_2567, net_2565, net_2563, net_2561, net_2559, net_2557, net_2555, net_2553, net_2568, net_2566, net_2564, net_2562, net_2560, net_2558, net_2556, net_2554}),
    .B({net_2361, net_2359, net_2357, net_2355, net_2353, net_2351, net_2349, net_2347, net_2362, net_2360, net_2358, net_2356, net_2354, net_2352, net_2350, net_2348}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({dangling_wire_0, net_2787, net_2786, net_2785, net_2784, net_2783, net_2782, net_2781, net_2579, net_2578, net_2577, net_2576, net_2575, net_2574, net_2573, net_2572, net_2369, net_2368, net_2367, net_2366, net_2365, net_2364, net_2371, net_2370, net_2165, net_2164, net_2163, net_2162, net_2161, net_2160, net_2159, net_2158})
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_0_15_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_3627, net_3625, net_3623, net_3621, net_3619, net_3617, net_3615, net_3613, net_3628, net_3626, net_3624, net_3622, net_3620, net_3618, net_3616, net_3614}),
    .B({net_3421, net_3419, net_3417, net_3415, net_3413, net_3411, net_3409, net_3407, net_3422, net_3420, net_3418, net_3416, net_3414, net_3412, net_3410, net_3408}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({dangling_wire_1, net_3847, net_3846, net_3845, net_3844, net_3843, net_3842, net_3841, net_3639, net_3638, net_3637, net_3636, net_3635, net_3634, net_3633, net_3632, net_3429, net_3428, net_3427, net_3426, net_3425, net_3424, net_3431, net_3430, net_3225, net_3224, net_3223, net_3222, net_3221, net_3220, net_3219, net_3218})
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_0_23_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_5368, net_5366, net_5364, net_5362, net_5360, net_5358, net_5356, net_5354, net_5369, net_5367, net_5365, net_5363, net_5361, net_5359, net_5357, net_5355}),
    .B({net_5162, net_5160, net_5158, net_5156, net_5154, net_5152, net_5150, net_5148, net_5163, net_5161, net_5159, net_5157, net_5155, net_5153, net_5151, net_5149}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({dangling_wire_2, net_5588, net_5587, net_5586, net_5585, net_5584, net_5583, net_5582, net_5380, net_5379, net_5378, net_5377, net_5376, net_5375, net_5374, net_5373, net_5170, net_5169, net_5168, net_5167, net_5166, net_5165, net_5172, net_5171, net_4966, net_4965, net_4964, net_4963, net_4962, net_4961, net_4960, net_4959})
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_0_5_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_1507, net_1505, net_1503, net_1501, net_1499, net_1497, net_1495, net_1493, net_1508, net_1506, net_1504, net_1502, net_1500, net_1498, net_1496, net_1494}),
    .B({net_1301, net_1299, net_1297, net_1295, net_1293, net_1291, net_1289, net_1287, net_1302, net_1300, net_1298, net_1296, net_1294, net_1292, net_1290, net_1288}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({dangling_wire_3, net_1727, net_1726, net_1725, net_1724, net_1723, net_1722, net_1721, net_1519, net_1518, net_1517, net_1516, net_1515, net_1514, net_1513, net_1512, net_1309, net_1308, net_1307, net_1306, net_1305, net_1304, net_1311, net_1310, net_1105, net_1104, net_1103, net_1102, net_1101, net_1100, net_1099, net_1098})
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_25_10_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_100347, net_100345, net_100343, net_100341, net_100339, net_100337, net_100335, net_100333, net_100348, net_100346, net_100344, net_100342, net_100340, net_100338, net_100336, net_100334}),
    .B({net_100197, net_100195, net_100193, net_100191, net_100189, net_100187, net_100185, net_100183, net_100198, net_100196, net_100194, net_100192, net_100190, net_100188, net_100186, net_100184}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({net_100511, net_100510, net_100509, net_100508, net_100507, net_100506, net_100505, net_100504, net_100359, net_100358, net_100357, net_100356, net_100355, net_100354, net_100353, net_100352, net_100205, net_100204, net_100203, net_100202, net_100201, net_100200, net_100207, net_100206, net_100057, net_100056, net_100055, net_100054, net_100053, net_100052, net_100051, net_100050})
  );
  SB_MAC16_MAS_U_16X16_BYPASS MAC16_25_5_0 (
    .ACCUMCI(),
    .ACCUMCO(),
    .ADDSUBBOT(gnd),
    .ADDSUBTOP(gnd),
    .AHOLD(gnd),
    .BHOLD(gnd),
    .CE(),
    .CHOLD(gnd),
    .CI(gnd),
    .CLK(),
    .DHOLD(gnd),
    .IRSTBOT(),
    .IRSTTOP(),
    .OHOLDBOT(gnd),
    .OHOLDTOP(gnd),
    .OLOADBOT(gnd),
    .OLOADTOP(gnd),
    .ORSTBOT(),
    .ORSTTOP(),
    .SIGNEXTIN(),
    .SIGNEXTOUT(),
    .A({net_99567, net_99565, net_99563, net_99561, net_99559, net_99557, net_99555, net_99553, net_99568, net_99566, net_99564, net_99562, net_99560, net_99558, net_99556, net_99554}),
    .B({net_99417, net_99415, net_99413, net_99411, net_99409, net_99407, net_99405, net_99403, net_99418, net_99416, net_99414, net_99412, net_99410, net_99408, net_99406, net_99404}),
    .C({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .D({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
    .O({net_99731, net_99730, net_99729, net_99728, net_99727, net_99726, net_99725, net_99724, net_99579, net_99578, net_99577, net_99576, net_99575, net_99574, net_99573, net_99572, net_99425, net_99424, net_99423, net_99422, net_99421, net_99420, net_99427, net_99426, net_99277, net_99276, net_99275, net_99274, net_99273, net_99272, net_99271, net_99270})
  );
  InMux inmux_0_11_2315_2359 (
    .I(net_2315),
    .O(net_2359)
  );
  InMux inmux_0_11_2322_2352 (
    .I(net_2322),
    .O(net_2352)
  );
  InMux inmux_0_11_2327_2349 (
    .I(net_2327),
    .O(net_2349)
  );
  InMux inmux_0_11_2330_2350 (
    .I(net_2330),
    .O(net_2350)
  );
  InMux inmux_0_11_2331_2356 (
    .I(net_2331),
    .O(net_2356)
  );
  InMux inmux_0_11_2332_2353 (
    .I(net_2332),
    .O(net_2353)
  );
  InMux inmux_0_11_2333_2360 (
    .I(net_2333),
    .O(net_2360)
  );
  InMux inmux_0_11_2334_2354 (
    .I(net_2334),
    .O(net_2354)
  );
  InMux inmux_0_11_2336_2358 (
    .I(net_2336),
    .O(net_2358)
  );
  InMux inmux_0_11_2337_2355 (
    .I(net_2337),
    .O(net_2355)
  );
  InMux inmux_0_11_2338_2351 (
    .I(net_2338),
    .O(net_2351)
  );
  InMux inmux_0_11_2339_2362 (
    .I(net_2339),
    .O(net_2362)
  );
  InMux inmux_0_11_2340_2348 (
    .I(net_2340),
    .O(net_2348)
  );
  InMux inmux_0_11_2342_2347 (
    .I(net_2342),
    .O(net_2347)
  );
  InMux inmux_0_11_2343_2361 (
    .I(net_2343),
    .O(net_2361)
  );
  InMux inmux_0_11_2345_2357 (
    .I(net_2345),
    .O(net_2357)
  );
  InMux inmux_0_12_2520_2559 (
    .I(net_2520),
    .O(net_2559)
  );
  InMux inmux_0_12_2521_2561 (
    .I(net_2521),
    .O(net_2561)
  );
  InMux inmux_0_12_2522_2555 (
    .I(net_2522),
    .O(net_2555)
  );
  InMux inmux_0_12_2523_2553 (
    .I(net_2523),
    .O(net_2553)
  );
  InMux inmux_0_12_2524_2564 (
    .I(net_2524),
    .O(net_2564)
  );
  InMux inmux_0_12_2526_2567 (
    .I(net_2526),
    .O(net_2567)
  );
  InMux inmux_0_12_2528_2566 (
    .I(net_2528),
    .O(net_2566)
  );
  InMux inmux_0_12_2529_2556 (
    .I(net_2529),
    .O(net_2556)
  );
  InMux inmux_0_12_2530_2562 (
    .I(net_2530),
    .O(net_2562)
  );
  InMux inmux_0_12_2531_2563 (
    .I(net_2531),
    .O(net_2563)
  );
  InMux inmux_0_12_2533_2568 (
    .I(net_2533),
    .O(net_2568)
  );
  InMux inmux_0_12_2534_2557 (
    .I(net_2534),
    .O(net_2557)
  );
  InMux inmux_0_12_2535_2560 (
    .I(net_2535),
    .O(net_2560)
  );
  InMux inmux_0_12_2544_2565 (
    .I(net_2544),
    .O(net_2565)
  );
  InMux inmux_0_12_2546_2558 (
    .I(net_2546),
    .O(net_2558)
  );
  InMux inmux_0_12_2548_2554 (
    .I(net_2548),
    .O(net_2554)
  );
  InMux inmux_0_16_3380_3410 (
    .I(net_3380),
    .O(net_3410)
  );
  InMux inmux_0_16_3382_3416 (
    .I(net_3382),
    .O(net_3416)
  );
  InMux inmux_0_16_3383_3414 (
    .I(net_3383),
    .O(net_3414)
  );
  InMux inmux_0_16_3385_3418 (
    .I(net_3385),
    .O(net_3418)
  );
  InMux inmux_0_16_3386_3411 (
    .I(net_3386),
    .O(net_3411)
  );
  InMux inmux_0_16_3388_3407 (
    .I(net_3388),
    .O(net_3407)
  );
  InMux inmux_0_16_3389_3422 (
    .I(net_3389),
    .O(net_3422)
  );
  InMux inmux_0_16_3390_3421 (
    .I(net_3390),
    .O(net_3421)
  );
  InMux inmux_0_16_3392_3417 (
    .I(net_3392),
    .O(net_3417)
  );
  InMux inmux_0_16_3393_3408 (
    .I(net_3393),
    .O(net_3408)
  );
  InMux inmux_0_16_3394_3409 (
    .I(net_3394),
    .O(net_3409)
  );
  InMux inmux_0_16_3395_3420 (
    .I(net_3395),
    .O(net_3420)
  );
  InMux inmux_0_16_3397_3412 (
    .I(net_3397),
    .O(net_3412)
  );
  InMux inmux_0_16_3399_3413 (
    .I(net_3399),
    .O(net_3413)
  );
  InMux inmux_0_16_3400_3419 (
    .I(net_3400),
    .O(net_3419)
  );
  InMux inmux_0_16_3402_3415 (
    .I(net_3402),
    .O(net_3415)
  );
  InMux inmux_0_17_3580_3615 (
    .I(net_3580),
    .O(net_3615)
  );
  InMux inmux_0_17_3582_3627 (
    .I(net_3582),
    .O(net_3627)
  );
  InMux inmux_0_17_3583_3626 (
    .I(net_3583),
    .O(net_3626)
  );
  InMux inmux_0_17_3585_3617 (
    .I(net_3585),
    .O(net_3617)
  );
  InMux inmux_0_17_3587_3625 (
    .I(net_3587),
    .O(net_3625)
  );
  InMux inmux_0_17_3589_3619 (
    .I(net_3589),
    .O(net_3619)
  );
  InMux inmux_0_17_3590_3621 (
    .I(net_3590),
    .O(net_3621)
  );
  InMux inmux_0_17_3592_3622 (
    .I(net_3592),
    .O(net_3622)
  );
  InMux inmux_0_17_3594_3613 (
    .I(net_3594),
    .O(net_3613)
  );
  InMux inmux_0_17_3595_3624 (
    .I(net_3595),
    .O(net_3624)
  );
  InMux inmux_0_17_3597_3614 (
    .I(net_3597),
    .O(net_3614)
  );
  InMux inmux_0_17_3598_3628 (
    .I(net_3598),
    .O(net_3628)
  );
  InMux inmux_0_17_3600_3616 (
    .I(net_3600),
    .O(net_3616)
  );
  InMux inmux_0_17_3606_3618 (
    .I(net_3606),
    .O(net_3618)
  );
  InMux inmux_0_17_3607_3623 (
    .I(net_3607),
    .O(net_3623)
  );
  InMux inmux_0_17_3611_3620 (
    .I(net_3611),
    .O(net_3620)
  );
  InMux inmux_0_24_5117_5151 (
    .I(net_5117),
    .O(net_5151)
  );
  InMux inmux_0_24_5118_5149 (
    .I(net_5118),
    .O(net_5149)
  );
  InMux inmux_0_24_5120_5160 (
    .I(net_5120),
    .O(net_5160)
  );
  InMux inmux_0_24_5122_5161 (
    .I(net_5122),
    .O(net_5161)
  );
  InMux inmux_0_24_5123_5157 (
    .I(net_5123),
    .O(net_5157)
  );
  InMux inmux_0_24_5125_5148 (
    .I(net_5125),
    .O(net_5148)
  );
  InMux inmux_0_24_5126_5163 (
    .I(net_5126),
    .O(net_5163)
  );
  InMux inmux_0_24_5127_5156 (
    .I(net_5127),
    .O(net_5156)
  );
  InMux inmux_0_24_5128_5150 (
    .I(net_5128),
    .O(net_5150)
  );
  InMux inmux_0_24_5133_5162 (
    .I(net_5133),
    .O(net_5162)
  );
  InMux inmux_0_24_5134_5152 (
    .I(net_5134),
    .O(net_5152)
  );
  InMux inmux_0_24_5140_5158 (
    .I(net_5140),
    .O(net_5158)
  );
  InMux inmux_0_24_5141_5153 (
    .I(net_5141),
    .O(net_5153)
  );
  InMux inmux_0_24_5142_5159 (
    .I(net_5142),
    .O(net_5159)
  );
  InMux inmux_0_24_5144_5155 (
    .I(net_5144),
    .O(net_5155)
  );
  InMux inmux_0_24_5146_5154 (
    .I(net_5146),
    .O(net_5154)
  );
  InMux inmux_0_25_5323_5365 (
    .I(net_5323),
    .O(net_5365)
  );
  InMux inmux_0_25_5325_5360 (
    .I(net_5325),
    .O(net_5360)
  );
  InMux inmux_0_25_5326_5354 (
    .I(net_5326),
    .O(net_5354)
  );
  InMux inmux_0_25_5327_5356 (
    .I(net_5327),
    .O(net_5356)
  );
  InMux inmux_0_25_5328_5362 (
    .I(net_5328),
    .O(net_5362)
  );
  InMux inmux_0_25_5329_5355 (
    .I(net_5329),
    .O(net_5355)
  );
  InMux inmux_0_25_5330_5369 (
    .I(net_5330),
    .O(net_5369)
  );
  InMux inmux_0_25_5331_5367 (
    .I(net_5331),
    .O(net_5367)
  );
  InMux inmux_0_25_5332_5364 (
    .I(net_5332),
    .O(net_5364)
  );
  InMux inmux_0_25_5336_5368 (
    .I(net_5336),
    .O(net_5368)
  );
  InMux inmux_0_25_5340_5366 (
    .I(net_5340),
    .O(net_5366)
  );
  InMux inmux_0_25_5341_5361 (
    .I(net_5341),
    .O(net_5361)
  );
  InMux inmux_0_25_5342_5358 (
    .I(net_5342),
    .O(net_5358)
  );
  InMux inmux_0_25_5344_5363 (
    .I(net_5344),
    .O(net_5363)
  );
  InMux inmux_0_25_5345_5359 (
    .I(net_5345),
    .O(net_5359)
  );
  InMux inmux_0_25_5346_5357 (
    .I(net_5346),
    .O(net_5357)
  );
  InMux inmux_0_6_1257_1296 (
    .I(net_1257),
    .O(net_1296)
  );
  InMux inmux_0_6_1258_1298 (
    .I(net_1258),
    .O(net_1298)
  );
  InMux inmux_0_6_1259_1300 (
    .I(net_1259),
    .O(net_1300)
  );
  InMux inmux_0_6_1262_1299 (
    .I(net_1262),
    .O(net_1299)
  );
  InMux inmux_0_6_1264_1295 (
    .I(net_1264),
    .O(net_1295)
  );
  InMux inmux_0_6_1267_1290 (
    .I(net_1267),
    .O(net_1290)
  );
  InMux inmux_0_6_1268_1287 (
    .I(net_1268),
    .O(net_1287)
  );
  InMux inmux_0_6_1272_1301 (
    .I(net_1272),
    .O(net_1301)
  );
  InMux inmux_0_6_1274_1293 (
    .I(net_1274),
    .O(net_1293)
  );
  InMux inmux_0_6_1275_1291 (
    .I(net_1275),
    .O(net_1291)
  );
  InMux inmux_0_6_1276_1302 (
    .I(net_1276),
    .O(net_1302)
  );
  InMux inmux_0_6_1278_1288 (
    .I(net_1278),
    .O(net_1288)
  );
  InMux inmux_0_6_1279_1294 (
    .I(net_1279),
    .O(net_1294)
  );
  InMux inmux_0_6_1280_1292 (
    .I(net_1280),
    .O(net_1292)
  );
  InMux inmux_0_6_1281_1297 (
    .I(net_1281),
    .O(net_1297)
  );
  InMux inmux_0_6_1285_1289 (
    .I(net_1285),
    .O(net_1289)
  );
  InMux inmux_0_7_1461_1501 (
    .I(net_1461),
    .O(net_1501)
  );
  InMux inmux_0_7_1464_1503 (
    .I(net_1464),
    .O(net_1503)
  );
  InMux inmux_0_7_1471_1496 (
    .I(net_1471),
    .O(net_1496)
  );
  InMux inmux_0_7_1474_1494 (
    .I(net_1474),
    .O(net_1494)
  );
  InMux inmux_0_7_1476_1508 (
    .I(net_1476),
    .O(net_1508)
  );
  InMux inmux_0_7_1478_1499 (
    .I(net_1478),
    .O(net_1499)
  );
  InMux inmux_0_7_1479_1497 (
    .I(net_1479),
    .O(net_1497)
  );
  InMux inmux_0_7_1483_1506 (
    .I(net_1483),
    .O(net_1506)
  );
  InMux inmux_0_7_1484_1505 (
    .I(net_1484),
    .O(net_1505)
  );
  InMux inmux_0_7_1485_1495 (
    .I(net_1485),
    .O(net_1495)
  );
  InMux inmux_0_7_1486_1498 (
    .I(net_1486),
    .O(net_1498)
  );
  InMux inmux_0_7_1487_1504 (
    .I(net_1487),
    .O(net_1504)
  );
  InMux inmux_0_7_1488_1502 (
    .I(net_1488),
    .O(net_1502)
  );
  InMux inmux_0_7_1489_1507 (
    .I(net_1489),
    .O(net_1507)
  );
  InMux inmux_0_7_1490_1493 (
    .I(net_1490),
    .O(net_1493)
  );
  InMux inmux_0_7_1491_1500 (
    .I(net_1491),
    .O(net_1500)
  );
  InMux inmux_10_10_42436_42500 (
    .I(net_42436),
    .O(net_42500)
  );
  InMux inmux_10_10_42437_42480 (
    .I(net_42437),
    .O(net_42480)
  );
  InMux inmux_10_10_42439_42506 (
    .I(net_42439),
    .O(net_42506)
  );
  InMux inmux_10_10_42444_42470 (
    .I(net_42444),
    .O(net_42470)
  );
  InMux inmux_10_10_42445_42512 (
    .I(net_42445),
    .O(net_42512)
  );
  InMux inmux_10_10_42448_42475 (
    .I(net_42448),
    .O(net_42475)
  );
  InMux inmux_10_10_42454_42505 (
    .I(net_42454),
    .O(net_42505)
  );
  InMux inmux_10_10_42456_42486 (
    .I(net_42456),
    .O(net_42486)
  );
  ClkMux inmux_10_10_5_42515 (
    .I(net_5),
    .O(net_42515)
  );
  SRMux inmux_10_10_9_42516 (
    .I(net_9),
    .O(net_42516)
  );
  InMux inmux_10_11_42558_42634 (
    .I(net_42558),
    .O(net_42634)
  );
  InMux inmux_10_11_42559_42616 (
    .I(net_42559),
    .O(net_42616)
  );
  InMux inmux_10_11_42560_42615 (
    .I(net_42560),
    .O(net_42615)
  );
  InMux inmux_10_11_42560_42636 (
    .I(net_42560),
    .O(net_42636)
  );
  InMux inmux_10_11_42565_42633 (
    .I(net_42565),
    .O(net_42633)
  );
  InMux inmux_10_11_42567_42598 (
    .I(net_42567),
    .O(net_42598)
  );
  InMux inmux_10_11_42569_42617 (
    .I(net_42569),
    .O(net_42617)
  );
  InMux inmux_10_11_42572_42609 (
    .I(net_42572),
    .O(net_42609)
  );
  InMux inmux_10_11_42575_42618 (
    .I(net_42575),
    .O(net_42618)
  );
  InMux inmux_10_11_42575_42635 (
    .I(net_42575),
    .O(net_42635)
  );
  CEMux inmux_10_11_42576_42637 (
    .I(net_42576),
    .O(net_42637)
  );
  InMux inmux_10_11_42581_42594 (
    .I(net_42581),
    .O(net_42594)
  );
  InMux inmux_10_11_42588_42630 (
    .I(net_42588),
    .O(net_42630)
  );
  ClkMux inmux_10_11_5_42638 (
    .I(net_5),
    .O(net_42638)
  );
  InMux inmux_10_12_42683_42726 (
    .I(net_42683),
    .O(net_42726)
  );
  CEMux inmux_10_12_42692_42760 (
    .I(net_42692),
    .O(net_42760)
  );
  ClkMux inmux_10_12_5_42761 (
    .I(net_5),
    .O(net_42761)
  );
  CEMux inmux_10_13_42806_42883 (
    .I(net_42806),
    .O(net_42883)
  );
  InMux inmux_10_13_42810_42851 (
    .I(net_42810),
    .O(net_42851)
  );
  InMux inmux_10_13_42814_42843 (
    .I(net_42814),
    .O(net_42843)
  );
  ClkMux inmux_10_13_5_42884 (
    .I(net_5),
    .O(net_42884)
  );
  InMux inmux_10_14_42927_43003 (
    .I(net_42927),
    .O(net_43003)
  );
  InMux inmux_10_14_42936_42969 (
    .I(net_42936),
    .O(net_42969)
  );
  InMux inmux_10_14_42951_42961 (
    .I(net_42951),
    .O(net_42961)
  );
  InMux inmux_10_14_42952_42993 (
    .I(net_42952),
    .O(net_42993)
  );
  InMux inmux_10_14_42953_42985 (
    .I(net_42953),
    .O(net_42985)
  );
  CEMux inmux_10_14_42954_43006 (
    .I(net_42954),
    .O(net_43006)
  );
  InMux inmux_10_14_42955_42980 (
    .I(net_42955),
    .O(net_42980)
  );
  ClkMux inmux_10_14_5_43007 (
    .I(net_5),
    .O(net_43007)
  );
  CEMux inmux_10_15_43052_43129 (
    .I(net_43052),
    .O(net_43129)
  );
  InMux inmux_10_15_43053_43098 (
    .I(net_43053),
    .O(net_43098)
  );
  InMux inmux_10_15_43056_43109 (
    .I(net_43056),
    .O(net_43109)
  );
  InMux inmux_10_15_43061_43085 (
    .I(net_43061),
    .O(net_43085)
  );
  InMux inmux_10_15_43063_43128 (
    .I(net_43063),
    .O(net_43128)
  );
  InMux inmux_10_15_43065_43097 (
    .I(net_43065),
    .O(net_43097)
  );
  InMux inmux_10_15_43076_43096 (
    .I(net_43076),
    .O(net_43096)
  );
  InMux inmux_10_15_43077_43095 (
    .I(net_43077),
    .O(net_43095)
  );
  ClkMux inmux_10_15_5_43130 (
    .I(net_5),
    .O(net_43130)
  );
  InMux inmux_10_16_43182_43215 (
    .I(net_43182),
    .O(net_43215)
  );
  InMux inmux_10_16_43187_43226 (
    .I(net_43187),
    .O(net_43226)
  );
  CEMux inmux_10_16_43191_43252 (
    .I(net_43191),
    .O(net_43252)
  );
  InMux inmux_10_16_43192_43231 (
    .I(net_43192),
    .O(net_43231)
  );
  InMux inmux_10_16_43193_43237 (
    .I(net_43193),
    .O(net_43237)
  );
  InMux inmux_10_16_43196_43207 (
    .I(net_43196),
    .O(net_43207)
  );
  ClkMux inmux_10_16_5_43253 (
    .I(net_5),
    .O(net_43253)
  );
  InMux inmux_10_17_43296_43343 (
    .I(net_43296),
    .O(net_43343)
  );
  CEMux inmux_10_17_43298_43375 (
    .I(net_43298),
    .O(net_43375)
  );
  InMux inmux_10_17_43299_43330 (
    .I(net_43299),
    .O(net_43330)
  );
  InMux inmux_10_17_43299_43344 (
    .I(net_43299),
    .O(net_43344)
  );
  InMux inmux_10_17_43299_43366 (
    .I(net_43299),
    .O(net_43366)
  );
  InMux inmux_10_17_43300_43367 (
    .I(net_43300),
    .O(net_43367)
  );
  InMux inmux_10_17_43301_43332 (
    .I(net_43301),
    .O(net_43332)
  );
  InMux inmux_10_17_43302_43353 (
    .I(net_43302),
    .O(net_43353)
  );
  InMux inmux_10_17_43305_43372 (
    .I(net_43305),
    .O(net_43372)
  );
  InMux inmux_10_17_43307_43331 (
    .I(net_43307),
    .O(net_43331)
  );
  InMux inmux_10_17_43307_43341 (
    .I(net_43307),
    .O(net_43341)
  );
  InMux inmux_10_17_43307_43365 (
    .I(net_43307),
    .O(net_43365)
  );
  InMux inmux_10_17_43310_43335 (
    .I(net_43310),
    .O(net_43335)
  );
  InMux inmux_10_17_43315_43368 (
    .I(net_43315),
    .O(net_43368)
  );
  InMux inmux_10_17_43316_43329 (
    .I(net_43316),
    .O(net_43329)
  );
  InMux inmux_10_17_43319_43342 (
    .I(net_43319),
    .O(net_43342)
  );
  ClkMux inmux_10_17_5_43376 (
    .I(net_5),
    .O(net_43376)
  );
  InMux inmux_10_18_43419_43454 (
    .I(net_43419),
    .O(net_43454)
  );
  InMux inmux_10_18_43421_43466 (
    .I(net_43421),
    .O(net_43466)
  );
  InMux inmux_10_18_43422_43460 (
    .I(net_43422),
    .O(net_43460)
  );
  InMux inmux_10_18_43425_43488 (
    .I(net_43425),
    .O(net_43488)
  );
  InMux inmux_10_18_43426_43467 (
    .I(net_43426),
    .O(net_43467)
  );
  InMux inmux_10_18_43428_43452 (
    .I(net_43428),
    .O(net_43452)
  );
  InMux inmux_10_18_43431_43453 (
    .I(net_43431),
    .O(net_43453)
  );
  InMux inmux_10_18_43431_43458 (
    .I(net_43431),
    .O(net_43458)
  );
  InMux inmux_10_18_43431_43465 (
    .I(net_43431),
    .O(net_43465)
  );
  InMux inmux_10_18_43431_43470 (
    .I(net_43431),
    .O(net_43470)
  );
  InMux inmux_10_18_43431_43477 (
    .I(net_43431),
    .O(net_43477)
  );
  InMux inmux_10_18_43431_43484 (
    .I(net_43431),
    .O(net_43484)
  );
  InMux inmux_10_18_43431_43489 (
    .I(net_43431),
    .O(net_43489)
  );
  InMux inmux_10_18_43431_43496 (
    .I(net_43431),
    .O(net_43496)
  );
  InMux inmux_10_18_43432_43495 (
    .I(net_43432),
    .O(net_43495)
  );
  InMux inmux_10_18_43434_43485 (
    .I(net_43434),
    .O(net_43485)
  );
  InMux inmux_10_18_43435_43473 (
    .I(net_43435),
    .O(net_43473)
  );
  InMux inmux_10_18_43437_43478 (
    .I(net_43437),
    .O(net_43478)
  );
  InMux inmux_10_18_43438_43491 (
    .I(net_43438),
    .O(net_43491)
  );
  InMux inmux_10_18_43439_43476 (
    .I(net_43439),
    .O(net_43476)
  );
  InMux inmux_10_18_43441_43459 (
    .I(net_43441),
    .O(net_43459)
  );
  InMux inmux_10_18_43444_43471 (
    .I(net_43444),
    .O(net_43471)
  );
  InMux inmux_10_18_43448_43497 (
    .I(net_43448),
    .O(net_43497)
  );
  InMux inmux_10_18_43450_43483 (
    .I(net_43450),
    .O(net_43483)
  );
  ClkMux inmux_10_18_5_43499 (
    .I(net_5),
    .O(net_43499)
  );
  CEMux inmux_10_18_6_43498 (
    .I(net_6),
    .O(net_43498)
  );
  SRMux inmux_10_18_9_43500 (
    .I(net_9),
    .O(net_43500)
  );
  CEMux inmux_10_19_43544_43621 (
    .I(net_43544),
    .O(net_43621)
  );
  InMux inmux_10_19_43549_43619 (
    .I(net_43549),
    .O(net_43619)
  );
  InMux inmux_10_19_43551_43584 (
    .I(net_43551),
    .O(net_43584)
  );
  InMux inmux_10_19_43551_43618 (
    .I(net_43551),
    .O(net_43618)
  );
  InMux inmux_10_19_43556_43617 (
    .I(net_43556),
    .O(net_43617)
  );
  InMux inmux_10_19_43557_43582 (
    .I(net_43557),
    .O(net_43582)
  );
  InMux inmux_10_19_43559_43581 (
    .I(net_43559),
    .O(net_43581)
  );
  InMux inmux_10_19_43568_43583 (
    .I(net_43568),
    .O(net_43583)
  );
  InMux inmux_10_19_43569_43620 (
    .I(net_43569),
    .O(net_43620)
  );
  ClkMux inmux_10_19_5_43622 (
    .I(net_5),
    .O(net_43622)
  );
  SRMux inmux_10_19_9_43623 (
    .I(net_9),
    .O(net_43623)
  );
  InMux inmux_10_1_41289_41358 (
    .I(net_41289),
    .O(net_41358)
  );
  InMux inmux_10_1_41292_41333 (
    .I(net_41292),
    .O(net_41333)
  );
  InMux inmux_10_1_41293_41329 (
    .I(net_41293),
    .O(net_41329)
  );
  InMux inmux_10_1_41294_41323 (
    .I(net_41294),
    .O(net_41323)
  );
  InMux inmux_10_1_41294_41366 (
    .I(net_41294),
    .O(net_41366)
  );
  InMux inmux_10_1_41299_41352 (
    .I(net_41299),
    .O(net_41352)
  );
  InMux inmux_10_1_41302_41334 (
    .I(net_41302),
    .O(net_41334)
  );
  InMux inmux_10_1_41303_41328 (
    .I(net_41303),
    .O(net_41328)
  );
  InMux inmux_10_1_41309_41322 (
    .I(net_41309),
    .O(net_41322)
  );
  InMux inmux_10_1_41309_41365 (
    .I(net_41309),
    .O(net_41365)
  );
  InMux inmux_10_1_41320_41330 (
    .I(net_41320),
    .O(net_41330)
  );
  InMux inmux_10_1_41326_41336 (
    .I(net_41326),
    .O(net_41336)
  );
  ClkMux inmux_10_1_5_41368 (
    .I(net_5),
    .O(net_41368)
  );
  SRMux inmux_10_1_9_41369 (
    .I(net_9),
    .O(net_41369)
  );
  InMux inmux_10_2_41452_41526 (
    .I(net_41452),
    .O(net_41526)
  );
  InMux inmux_10_2_41457_41517 (
    .I(net_41457),
    .O(net_41517)
  );
  InMux inmux_10_2_41458_41504 (
    .I(net_41458),
    .O(net_41504)
  );
  InMux inmux_10_2_41470_41511 (
    .I(net_41470),
    .O(net_41511)
  );
  InMux inmux_10_2_41474_41521 (
    .I(net_41474),
    .O(net_41521)
  );
  InMux inmux_10_2_41475_41497 (
    .I(net_41475),
    .O(net_41497)
  );
  InMux inmux_10_2_41477_41490 (
    .I(net_41477),
    .O(net_41490)
  );
  InMux inmux_10_2_41479_41485 (
    .I(net_41479),
    .O(net_41485)
  );
  ClkMux inmux_10_2_5_41531 (
    .I(net_5),
    .O(net_41531)
  );
  SRMux inmux_10_2_9_41532 (
    .I(net_9),
    .O(net_41532)
  );
  InMux inmux_10_3_41584_41637 (
    .I(net_41584),
    .O(net_41637)
  );
  InMux inmux_10_3_41589_41633 (
    .I(net_41589),
    .O(net_41633)
  );
  InMux inmux_10_3_41593_41615 (
    .I(net_41593),
    .O(net_41615)
  );
  InMux inmux_10_3_41594_41650 (
    .I(net_41594),
    .O(net_41650)
  );
  InMux inmux_10_3_41595_41608 (
    .I(net_41595),
    .O(net_41608)
  );
  InMux inmux_10_3_41598_41622 (
    .I(net_41598),
    .O(net_41622)
  );
  InMux inmux_10_3_41603_41645 (
    .I(net_41603),
    .O(net_41645)
  );
  InMux inmux_10_3_41604_41627 (
    .I(net_41604),
    .O(net_41627)
  );
  ClkMux inmux_10_3_5_41654 (
    .I(net_5),
    .O(net_41654)
  );
  SRMux inmux_10_3_9_41655 (
    .I(net_9),
    .O(net_41655)
  );
  InMux inmux_10_4_41703_41730 (
    .I(net_41703),
    .O(net_41730)
  );
  InMux inmux_10_4_41704_41750 (
    .I(net_41704),
    .O(net_41750)
  );
  InMux inmux_10_4_41706_41737 (
    .I(net_41706),
    .O(net_41737)
  );
  InMux inmux_10_4_41708_41732 (
    .I(net_41708),
    .O(net_41732)
  );
  InMux inmux_10_4_41710_41775 (
    .I(net_41710),
    .O(net_41775)
  );
  InMux inmux_10_4_41712_41773 (
    .I(net_41712),
    .O(net_41773)
  );
  InMux inmux_10_4_41714_41731 (
    .I(net_41714),
    .O(net_41731)
  );
  InMux inmux_10_4_41719_41761 (
    .I(net_41719),
    .O(net_41761)
  );
  InMux inmux_10_4_41724_41766 (
    .I(net_41724),
    .O(net_41766)
  );
  InMux inmux_10_4_41725_41733 (
    .I(net_41725),
    .O(net_41733)
  );
  InMux inmux_10_4_41725_41772 (
    .I(net_41725),
    .O(net_41772)
  );
  InMux inmux_10_4_41727_41774 (
    .I(net_41727),
    .O(net_41774)
  );
  ClkMux inmux_10_4_5_41777 (
    .I(net_5),
    .O(net_41777)
  );
  CEMux inmux_10_4_8_41776 (
    .I(net_8),
    .O(net_41776)
  );
  InMux inmux_10_5_41828_41859 (
    .I(net_41828),
    .O(net_41859)
  );
  InMux inmux_10_5_41832_41895 (
    .I(net_41832),
    .O(net_41895)
  );
  InMux inmux_10_5_41842_41886 (
    .I(net_41842),
    .O(net_41886)
  );
  InMux inmux_10_5_41846_41892 (
    .I(net_41846),
    .O(net_41892)
  );
  InMux inmux_10_5_41849_41877 (
    .I(net_41849),
    .O(net_41877)
  );
  ClkMux inmux_10_5_5_41900 (
    .I(net_5),
    .O(net_41900)
  );
  SRMux inmux_10_5_9_41901 (
    .I(net_9),
    .O(net_41901)
  );
  CEMux inmux_10_6_10_42022 (
    .I(net_10),
    .O(net_42022)
  );
  InMux inmux_10_6_41953_42001 (
    .I(net_41953),
    .O(net_42001)
  );
  InMux inmux_10_6_41960_42018 (
    .I(net_41960),
    .O(net_42018)
  );
  InMux inmux_10_6_41968_41983 (
    .I(net_41968),
    .O(net_41983)
  );
  ClkMux inmux_10_6_5_42023 (
    .I(net_5),
    .O(net_42023)
  );
  InMux inmux_10_7_42070_42144 (
    .I(net_42070),
    .O(net_42144)
  );
  InMux inmux_10_7_42072_42125 (
    .I(net_42072),
    .O(net_42125)
  );
  InMux inmux_10_7_42073_42100 (
    .I(net_42073),
    .O(net_42100)
  );
  InMux inmux_10_7_42074_42107 (
    .I(net_42074),
    .O(net_42107)
  );
  InMux inmux_10_7_42082_42123 (
    .I(net_42082),
    .O(net_42123)
  );
  InMux inmux_10_7_42091_42130 (
    .I(net_42091),
    .O(net_42130)
  );
  InMux inmux_10_7_42093_42118 (
    .I(net_42093),
    .O(net_42118)
  );
  ClkMux inmux_10_7_5_42146 (
    .I(net_5),
    .O(net_42146)
  );
  SRMux inmux_10_7_9_42147 (
    .I(net_9),
    .O(net_42147)
  );
  InMux inmux_10_8_42193_42248 (
    .I(net_42193),
    .O(net_42248)
  );
  InMux inmux_10_8_42198_42255 (
    .I(net_42198),
    .O(net_42255)
  );
  InMux inmux_10_8_42199_42259 (
    .I(net_42199),
    .O(net_42259)
  );
  InMux inmux_10_8_42202_42229 (
    .I(net_42202),
    .O(net_42229)
  );
  InMux inmux_10_8_42203_42240 (
    .I(net_42203),
    .O(net_42240)
  );
  InMux inmux_10_8_42213_42225 (
    .I(net_42213),
    .O(net_42225)
  );
  InMux inmux_10_8_42218_42265 (
    .I(net_42218),
    .O(net_42265)
  );
  ClkMux inmux_10_8_5_42269 (
    .I(net_5),
    .O(net_42269)
  );
  SRMux inmux_10_8_9_42270 (
    .I(net_9),
    .O(net_42270)
  );
  CEMux inmux_10_9_10_42391 (
    .I(net_10),
    .O(net_42391)
  );
  InMux inmux_10_9_42319_42365 (
    .I(net_42319),
    .O(net_42365)
  );
  ClkMux inmux_10_9_5_42392 (
    .I(net_5),
    .O(net_42392)
  );
  CEMux inmux_11_10_46268_46345 (
    .I(net_46268),
    .O(net_46345)
  );
  InMux inmux_11_10_46273_46307 (
    .I(net_46273),
    .O(net_46307)
  );
  InMux inmux_11_10_46283_46343 (
    .I(net_46283),
    .O(net_46343)
  );
  InMux inmux_11_10_46285_46324 (
    .I(net_46285),
    .O(net_46324)
  );
  ClkMux inmux_11_10_5_46346 (
    .I(net_5),
    .O(net_46346)
  );
  InMux inmux_11_11_46389_46429 (
    .I(net_46389),
    .O(net_46429)
  );
  InMux inmux_11_11_46392_46459 (
    .I(net_46392),
    .O(net_46459)
  );
  InMux inmux_11_11_46395_46424 (
    .I(net_46395),
    .O(net_46424)
  );
  InMux inmux_11_11_46397_46437 (
    .I(net_46397),
    .O(net_46437)
  );
  InMux inmux_11_11_46401_46425 (
    .I(net_46401),
    .O(net_46425)
  );
  InMux inmux_11_11_46402_46434 (
    .I(net_46402),
    .O(net_46434)
  );
  InMux inmux_11_11_46402_46443 (
    .I(net_46402),
    .O(net_46443)
  );
  InMux inmux_11_11_46402_46465 (
    .I(net_46402),
    .O(net_46465)
  );
  InMux inmux_11_11_46403_46447 (
    .I(net_46403),
    .O(net_46447)
  );
  InMux inmux_11_11_46405_46422 (
    .I(net_46405),
    .O(net_46422)
  );
  InMux inmux_11_11_46409_46455 (
    .I(net_46409),
    .O(net_46455)
  );
  InMux inmux_11_11_46410_46442 (
    .I(net_46410),
    .O(net_46442)
  );
  InMux inmux_11_11_46414_46467 (
    .I(net_46414),
    .O(net_46467)
  );
  InMux inmux_11_11_46417_46423 (
    .I(net_46417),
    .O(net_46423)
  );
  ClkMux inmux_11_11_5_46469 (
    .I(net_5),
    .O(net_46469)
  );
  SRMux inmux_11_11_9_46470 (
    .I(net_9),
    .O(net_46470)
  );
  InMux inmux_11_12_46512_46557 (
    .I(net_46512),
    .O(net_46557)
  );
  InMux inmux_11_12_46518_46552 (
    .I(net_46518),
    .O(net_46552)
  );
  InMux inmux_11_12_46519_46546 (
    .I(net_46519),
    .O(net_46546)
  );
  InMux inmux_11_12_46522_46577 (
    .I(net_46522),
    .O(net_46577)
  );
  InMux inmux_11_12_46523_46547 (
    .I(net_46523),
    .O(net_46547)
  );
  InMux inmux_11_12_46527_46571 (
    .I(net_46527),
    .O(net_46571)
  );
  InMux inmux_11_12_46529_46572 (
    .I(net_46529),
    .O(net_46572)
  );
  InMux inmux_11_12_46530_46569 (
    .I(net_46530),
    .O(net_46569)
  );
  InMux inmux_11_12_46535_46560 (
    .I(net_46535),
    .O(net_46560)
  );
  InMux inmux_11_12_46536_46570 (
    .I(net_46536),
    .O(net_46570)
  );
  InMux inmux_11_12_46538_46548 (
    .I(net_46538),
    .O(net_46548)
  );
  InMux inmux_11_12_46538_46551 (
    .I(net_46538),
    .O(net_46551)
  );
  InMux inmux_11_12_46538_46558 (
    .I(net_46538),
    .O(net_46558)
  );
  InMux inmux_11_12_46538_46575 (
    .I(net_46538),
    .O(net_46575)
  );
  InMux inmux_11_12_46540_46553 (
    .I(net_46540),
    .O(net_46553)
  );
  InMux inmux_11_12_46543_46576 (
    .I(net_46543),
    .O(net_46576)
  );
  ClkMux inmux_11_12_5_46592 (
    .I(net_5),
    .O(net_46592)
  );
  CEMux inmux_11_12_6_46591 (
    .I(net_6),
    .O(net_46591)
  );
  SRMux inmux_11_12_9_46593 (
    .I(net_9),
    .O(net_46593)
  );
  InMux inmux_11_13_46636_46681 (
    .I(net_46636),
    .O(net_46681)
  );
  InMux inmux_11_13_46644_46694 (
    .I(net_46644),
    .O(net_46694)
  );
  CEMux inmux_11_13_46653_46714 (
    .I(net_46653),
    .O(net_46714)
  );
  InMux inmux_11_13_46655_46680 (
    .I(net_46655),
    .O(net_46680)
  );
  InMux inmux_11_13_46660_46682 (
    .I(net_46660),
    .O(net_46682)
  );
  InMux inmux_11_13_46661_46683 (
    .I(net_46661),
    .O(net_46683)
  );
  ClkMux inmux_11_13_5_46715 (
    .I(net_5),
    .O(net_46715)
  );
  InMux inmux_11_14_46758_46834 (
    .I(net_46758),
    .O(net_46834)
  );
  InMux inmux_11_14_46761_46806 (
    .I(net_46761),
    .O(net_46806)
  );
  InMux inmux_11_14_46762_46824 (
    .I(net_46762),
    .O(net_46824)
  );
  InMux inmux_11_14_46768_46794 (
    .I(net_46768),
    .O(net_46794)
  );
  InMux inmux_11_14_46771_46817 (
    .I(net_46771),
    .O(net_46817)
  );
  CEMux inmux_11_14_46785_46837 (
    .I(net_46785),
    .O(net_46837)
  );
  ClkMux inmux_11_14_5_46838 (
    .I(net_5),
    .O(net_46838)
  );
  InMux inmux_11_15_46882_46958 (
    .I(net_46882),
    .O(net_46958)
  );
  InMux inmux_11_15_46885_46923 (
    .I(net_46885),
    .O(net_46923)
  );
  InMux inmux_11_15_46887_46959 (
    .I(net_46887),
    .O(net_46959)
  );
  InMux inmux_11_15_46896_46950 (
    .I(net_46896),
    .O(net_46950)
  );
  InMux inmux_11_15_46897_46928 (
    .I(net_46897),
    .O(net_46928)
  );
  CEMux inmux_11_15_46899_46960 (
    .I(net_46899),
    .O(net_46960)
  );
  InMux inmux_11_15_46901_46926 (
    .I(net_46901),
    .O(net_46926)
  );
  InMux inmux_11_15_46901_46957 (
    .I(net_46901),
    .O(net_46957)
  );
  InMux inmux_11_15_46902_46915 (
    .I(net_46902),
    .O(net_46915)
  );
  InMux inmux_11_15_46904_46929 (
    .I(net_46904),
    .O(net_46929)
  );
  InMux inmux_11_15_46910_46938 (
    .I(net_46910),
    .O(net_46938)
  );
  InMux inmux_11_15_46911_46927 (
    .I(net_46911),
    .O(net_46927)
  );
  InMux inmux_11_15_46911_46956 (
    .I(net_46911),
    .O(net_46956)
  );
  ClkMux inmux_11_15_5_46961 (
    .I(net_5),
    .O(net_46961)
  );
  InMux inmux_11_16_47008_47037 (
    .I(net_47008),
    .O(net_47037)
  );
  InMux inmux_11_16_47012_47055 (
    .I(net_47012),
    .O(net_47055)
  );
  InMux inmux_11_16_47013_47046 (
    .I(net_47013),
    .O(net_47046)
  );
  InMux inmux_11_16_47018_47038 (
    .I(net_47018),
    .O(net_47038)
  );
  InMux inmux_11_16_47018_47043 (
    .I(net_47018),
    .O(net_47043)
  );
  InMux inmux_11_16_47018_47057 (
    .I(net_47018),
    .O(net_47057)
  );
  InMux inmux_11_16_47018_47064 (
    .I(net_47018),
    .O(net_47064)
  );
  InMux inmux_11_16_47022_47056 (
    .I(net_47022),
    .O(net_47056)
  );
  InMux inmux_11_16_47023_47062 (
    .I(net_47023),
    .O(net_47062)
  );
  InMux inmux_11_16_47030_47045 (
    .I(net_47030),
    .O(net_47045)
  );
  InMux inmux_11_16_47031_47063 (
    .I(net_47031),
    .O(net_47063)
  );
  InMux inmux_11_16_47033_47039 (
    .I(net_47033),
    .O(net_47039)
  );
  ClkMux inmux_11_16_5_47084 (
    .I(net_5),
    .O(net_47084)
  );
  CEMux inmux_11_16_6_47083 (
    .I(net_6),
    .O(net_47083)
  );
  SRMux inmux_11_16_9_47085 (
    .I(net_9),
    .O(net_47085)
  );
  InMux inmux_11_17_47128_47185 (
    .I(net_47128),
    .O(net_47185)
  );
  InMux inmux_11_17_47129_47198 (
    .I(net_47129),
    .O(net_47198)
  );
  InMux inmux_11_17_47131_47205 (
    .I(net_47131),
    .O(net_47205)
  );
  InMux inmux_11_17_47132_47173 (
    .I(net_47132),
    .O(net_47173)
  );
  InMux inmux_11_17_47135_47190 (
    .I(net_47135),
    .O(net_47190)
  );
  InMux inmux_11_17_47136_47162 (
    .I(net_47136),
    .O(net_47162)
  );
  InMux inmux_11_17_47137_47199 (
    .I(net_47137),
    .O(net_47199)
  );
  InMux inmux_11_17_47138_47191 (
    .I(net_47138),
    .O(net_47191)
  );
  InMux inmux_11_17_47138_47196 (
    .I(net_47138),
    .O(net_47196)
  );
  InMux inmux_11_17_47141_47192 (
    .I(net_47141),
    .O(net_47192)
  );
  InMux inmux_11_17_47141_47197 (
    .I(net_47141),
    .O(net_47197)
  );
  InMux inmux_11_17_47143_47193 (
    .I(net_47143),
    .O(net_47193)
  );
  CEMux inmux_11_17_47145_47206 (
    .I(net_47145),
    .O(net_47206)
  );
  InMux inmux_11_17_47156_47181 (
    .I(net_47156),
    .O(net_47181)
  );
  ClkMux inmux_11_17_5_47207 (
    .I(net_5),
    .O(net_47207)
  );
  InMux inmux_11_18_47250_47314 (
    .I(net_47250),
    .O(net_47314)
  );
  InMux inmux_11_18_47251_47296 (
    .I(net_47251),
    .O(net_47296)
  );
  CEMux inmux_11_18_47252_47329 (
    .I(net_47252),
    .O(net_47329)
  );
  InMux inmux_11_18_47255_47291 (
    .I(net_47255),
    .O(net_47291)
  );
  InMux inmux_11_18_47256_47316 (
    .I(net_47256),
    .O(net_47316)
  );
  InMux inmux_11_18_47257_47289 (
    .I(net_47257),
    .O(net_47289)
  );
  InMux inmux_11_18_47257_47315 (
    .I(net_47257),
    .O(net_47315)
  );
  InMux inmux_11_18_47260_47313 (
    .I(net_47260),
    .O(net_47313)
  );
  InMux inmux_11_18_47263_47297 (
    .I(net_47263),
    .O(net_47297)
  );
  InMux inmux_11_18_47264_47325 (
    .I(net_47264),
    .O(net_47325)
  );
  InMux inmux_11_18_47265_47295 (
    .I(net_47265),
    .O(net_47295)
  );
  InMux inmux_11_18_47265_47326 (
    .I(net_47265),
    .O(net_47326)
  );
  InMux inmux_11_18_47266_47328 (
    .I(net_47266),
    .O(net_47328)
  );
  InMux inmux_11_18_47268_47290 (
    .I(net_47268),
    .O(net_47290)
  );
  InMux inmux_11_18_47277_47292 (
    .I(net_47277),
    .O(net_47292)
  );
  InMux inmux_11_18_47278_47327 (
    .I(net_47278),
    .O(net_47327)
  );
  InMux inmux_11_18_47280_47298 (
    .I(net_47280),
    .O(net_47298)
  );
  ClkMux inmux_11_18_5_47330 (
    .I(net_5),
    .O(net_47330)
  );
  CEMux inmux_11_19_12_47452 (
    .I(net_12),
    .O(net_47452)
  );
  InMux inmux_11_19_47382_47413 (
    .I(net_47382),
    .O(net_47413)
  );
  ClkMux inmux_11_19_5_47453 (
    .I(net_5),
    .O(net_47453)
  );
  InMux inmux_11_1_45135_45178 (
    .I(net_45135),
    .O(net_45178)
  );
  ClkMux inmux_11_1_5_45199 (
    .I(net_5),
    .O(net_45199)
  );
  SRMux inmux_11_1_9_45200 (
    .I(net_9),
    .O(net_45200)
  );
  InMux inmux_11_2_45283_45340 (
    .I(net_45283),
    .O(net_45340)
  );
  InMux inmux_11_2_45296_45357 (
    .I(net_45296),
    .O(net_45357)
  );
  InMux inmux_11_2_45299_45323 (
    .I(net_45299),
    .O(net_45323)
  );
  InMux inmux_11_2_45300_45353 (
    .I(net_45300),
    .O(net_45353)
  );
  InMux inmux_11_2_45301_45347 (
    .I(net_45301),
    .O(net_45347)
  );
  InMux inmux_11_2_45304_45317 (
    .I(net_45304),
    .O(net_45317)
  );
  InMux inmux_11_2_45305_45316 (
    .I(net_45305),
    .O(net_45316)
  );
  InMux inmux_11_2_45308_45328 (
    .I(net_45308),
    .O(net_45328)
  );
  InMux inmux_11_2_45311_45322 (
    .I(net_45311),
    .O(net_45322)
  );
  InMux inmux_11_2_45312_45345 (
    .I(net_45312),
    .O(net_45345)
  );
  InMux inmux_11_2_45313_45329 (
    .I(net_45313),
    .O(net_45329)
  );
  InMux inmux_11_2_45314_45324 (
    .I(net_45314),
    .O(net_45324)
  );
  InMux inmux_11_2_45320_45330 (
    .I(net_45320),
    .O(net_45330)
  );
  ClkMux inmux_11_2_5_45362 (
    .I(net_5),
    .O(net_45362)
  );
  SRMux inmux_11_2_9_45363 (
    .I(net_9),
    .O(net_45363)
  );
  InMux inmux_11_3_45408_45458 (
    .I(net_45408),
    .O(net_45458)
  );
  InMux inmux_11_3_45411_45440 (
    .I(net_45411),
    .O(net_45440)
  );
  InMux inmux_11_3_45412_45463 (
    .I(net_45412),
    .O(net_45463)
  );
  InMux inmux_11_3_45413_45475 (
    .I(net_45413),
    .O(net_45475)
  );
  InMux inmux_11_3_45414_45464 (
    .I(net_45414),
    .O(net_45464)
  );
  InMux inmux_11_3_45415_45446 (
    .I(net_45415),
    .O(net_45446)
  );
  InMux inmux_11_3_45417_45451 (
    .I(net_45417),
    .O(net_45451)
  );
  InMux inmux_11_3_45418_45476 (
    .I(net_45418),
    .O(net_45476)
  );
  InMux inmux_11_3_45420_45452 (
    .I(net_45420),
    .O(net_45452)
  );
  InMux inmux_11_3_45425_45469 (
    .I(net_45425),
    .O(net_45469)
  );
  InMux inmux_11_3_45427_45457 (
    .I(net_45427),
    .O(net_45457)
  );
  InMux inmux_11_3_45429_45470 (
    .I(net_45429),
    .O(net_45470)
  );
  InMux inmux_11_3_45430_45445 (
    .I(net_45430),
    .O(net_45445)
  );
  InMux inmux_11_3_45435_45439 (
    .I(net_45435),
    .O(net_45439)
  );
  InMux inmux_11_3_45437_45447 (
    .I(net_45437),
    .O(net_45447)
  );
  InMux inmux_11_3_45443_45453 (
    .I(net_45443),
    .O(net_45453)
  );
  InMux inmux_11_3_45449_45459 (
    .I(net_45449),
    .O(net_45459)
  );
  InMux inmux_11_3_45455_45465 (
    .I(net_45455),
    .O(net_45465)
  );
  InMux inmux_11_3_45461_45471 (
    .I(net_45461),
    .O(net_45471)
  );
  InMux inmux_11_3_45467_45477 (
    .I(net_45467),
    .O(net_45477)
  );
  InMux inmux_11_3_45473_45483 (
    .I(net_45473),
    .O(net_45483)
  );
  InMux inmux_11_4_45529_45569 (
    .I(net_45529),
    .O(net_45569)
  );
  InMux inmux_11_4_45532_45587 (
    .I(net_45532),
    .O(net_45587)
  );
  InMux inmux_11_4_45533_45562 (
    .I(net_45533),
    .O(net_45562)
  );
  InMux inmux_11_4_45534_45568 (
    .I(net_45534),
    .O(net_45568)
  );
  InMux inmux_11_4_45538_45574 (
    .I(net_45538),
    .O(net_45574)
  );
  InMux inmux_11_4_45539_45580 (
    .I(net_45539),
    .O(net_45580)
  );
  InMux inmux_11_4_45541_45592 (
    .I(net_45541),
    .O(net_45592)
  );
  InMux inmux_11_4_45542_45598 (
    .I(net_45542),
    .O(net_45598)
  );
  InMux inmux_11_4_45543_45604 (
    .I(net_45543),
    .O(net_45604)
  );
  InMux inmux_11_4_45546_45575 (
    .I(net_45546),
    .O(net_45575)
  );
  InMux inmux_11_4_45546_45599 (
    .I(net_45546),
    .O(net_45599)
  );
  InMux inmux_11_4_45554_45581 (
    .I(net_45554),
    .O(net_45581)
  );
  InMux inmux_11_4_45554_45586 (
    .I(net_45554),
    .O(net_45586)
  );
  InMux inmux_11_4_45554_45593 (
    .I(net_45554),
    .O(net_45593)
  );
  InMux inmux_11_4_45554_45605 (
    .I(net_45554),
    .O(net_45605)
  );
  InMux inmux_11_4_45557_45563 (
    .I(net_45557),
    .O(net_45563)
  );
  InMux inmux_11_4_45560_45570 (
    .I(net_45560),
    .O(net_45570)
  );
  InMux inmux_11_4_45566_45576 (
    .I(net_45566),
    .O(net_45576)
  );
  InMux inmux_11_4_45572_45582 (
    .I(net_45572),
    .O(net_45582)
  );
  InMux inmux_11_4_45578_45588 (
    .I(net_45578),
    .O(net_45588)
  );
  InMux inmux_11_4_45584_45594 (
    .I(net_45584),
    .O(net_45594)
  );
  InMux inmux_11_4_45590_45600 (
    .I(net_45590),
    .O(net_45600)
  );
  InMux inmux_11_4_45596_45606 (
    .I(net_45596),
    .O(net_45606)
  );
  ClkMux inmux_11_4_5_45608 (
    .I(net_5),
    .O(net_45608)
  );
  SRMux inmux_11_4_9_45609 (
    .I(net_9),
    .O(net_45609)
  );
  InMux inmux_11_5_45646_45687 (
    .I(net_45646),
    .O(net_45687)
  );
  InMux inmux_11_5_45653_45715 (
    .I(net_45653),
    .O(net_45715)
  );
  InMux inmux_11_5_45654_45685 (
    .I(net_45654),
    .O(net_45685)
  );
  InMux inmux_11_5_45654_45692 (
    .I(net_45654),
    .O(net_45692)
  );
  InMux inmux_11_5_45658_45711 (
    .I(net_45658),
    .O(net_45711)
  );
  InMux inmux_11_5_45662_45720 (
    .I(net_45662),
    .O(net_45720)
  );
  InMux inmux_11_5_45663_45702 (
    .I(net_45663),
    .O(net_45702)
  );
  InMux inmux_11_5_45665_45697 (
    .I(net_45665),
    .O(net_45697)
  );
  InMux inmux_11_5_45666_45727 (
    .I(net_45666),
    .O(net_45727)
  );
  InMux inmux_11_5_45683_45693 (
    .I(net_45683),
    .O(net_45693)
  );
  ClkMux inmux_11_5_5_45731 (
    .I(net_5),
    .O(net_45731)
  );
  SRMux inmux_11_5_9_45732 (
    .I(net_9),
    .O(net_45732)
  );
  InMux inmux_11_6_45790_45814 (
    .I(net_45790),
    .O(net_45814)
  );
  InMux inmux_11_6_45791_45834 (
    .I(net_45791),
    .O(net_45834)
  );
  InMux inmux_11_6_45793_45810 (
    .I(net_45793),
    .O(net_45810)
  );
  InMux inmux_11_6_45796_45850 (
    .I(net_45796),
    .O(net_45850)
  );
  ClkMux inmux_11_6_5_45854 (
    .I(net_5),
    .O(net_45854)
  );
  SRMux inmux_11_6_9_45855 (
    .I(net_9),
    .O(net_45855)
  );
  CEMux inmux_11_7_10_45976 (
    .I(net_10),
    .O(net_45976)
  );
  InMux inmux_11_7_45905_45960 (
    .I(net_45905),
    .O(net_45960)
  );
  InMux inmux_11_7_45909_45933 (
    .I(net_45909),
    .O(net_45933)
  );
  InMux inmux_11_7_45923_45957 (
    .I(net_45923),
    .O(net_45957)
  );
  ClkMux inmux_11_7_5_45977 (
    .I(net_5),
    .O(net_45977)
  );
  InMux inmux_11_8_46021_46066 (
    .I(net_46021),
    .O(net_46066)
  );
  InMux inmux_11_8_46025_46092 (
    .I(net_46025),
    .O(net_46092)
  );
  InMux inmux_11_8_46028_46095 (
    .I(net_46028),
    .O(net_46095)
  );
  InMux inmux_11_8_46031_46079 (
    .I(net_46031),
    .O(net_46079)
  );
  InMux inmux_11_8_46033_46084 (
    .I(net_46033),
    .O(net_46084)
  );
  InMux inmux_11_8_46034_46061 (
    .I(net_46034),
    .O(net_46061)
  );
  InMux inmux_11_8_46040_46055 (
    .I(net_46040),
    .O(net_46055)
  );
  InMux inmux_11_8_46042_46072 (
    .I(net_46042),
    .O(net_46072)
  );
  InMux inmux_11_8_46042_46086 (
    .I(net_46042),
    .O(net_46086)
  );
  InMux inmux_11_8_46042_46089 (
    .I(net_46042),
    .O(net_46089)
  );
  InMux inmux_11_8_46042_46096 (
    .I(net_46042),
    .O(net_46096)
  );
  InMux inmux_11_8_46043_46071 (
    .I(net_46043),
    .O(net_46071)
  );
  ClkMux inmux_11_8_5_46100 (
    .I(net_5),
    .O(net_46100)
  );
  SRMux inmux_11_8_9_46101 (
    .I(net_9),
    .O(net_46101)
  );
  InMux inmux_11_9_46144_46201 (
    .I(net_46144),
    .O(net_46201)
  );
  InMux inmux_11_9_46154_46221 (
    .I(net_46154),
    .O(net_46221)
  );
  InMux inmux_11_9_46158_46183 (
    .I(net_46158),
    .O(net_46183)
  );
  ClkMux inmux_11_9_5_46223 (
    .I(net_5),
    .O(net_46223)
  );
  SRMux inmux_11_9_9_46224 (
    .I(net_9),
    .O(net_46224)
  );
  InMux inmux_12_10_50097_50149 (
    .I(net_50097),
    .O(net_50149)
  );
  InMux inmux_12_10_50097_50168 (
    .I(net_50097),
    .O(net_50168)
  );
  InMux inmux_12_10_50100_50174 (
    .I(net_50100),
    .O(net_50174)
  );
  InMux inmux_12_10_50101_50166 (
    .I(net_50101),
    .O(net_50166)
  );
  InMux inmux_12_10_50108_50139 (
    .I(net_50108),
    .O(net_50139)
  );
  InMux inmux_12_10_50110_50154 (
    .I(net_50110),
    .O(net_50154)
  );
  InMux inmux_12_10_50122_50151 (
    .I(net_50122),
    .O(net_50151)
  );
  ClkMux inmux_12_10_5_50177 (
    .I(net_5),
    .O(net_50177)
  );
  SRMux inmux_12_10_9_50178 (
    .I(net_9),
    .O(net_50178)
  );
  InMux inmux_12_11_50222_50274 (
    .I(net_50222),
    .O(net_50274)
  );
  InMux inmux_12_11_50224_50291 (
    .I(net_50224),
    .O(net_50291)
  );
  InMux inmux_12_11_50227_50285 (
    .I(net_50227),
    .O(net_50285)
  );
  CEMux inmux_12_11_50231_50299 (
    .I(net_50231),
    .O(net_50299)
  );
  InMux inmux_12_11_50233_50265 (
    .I(net_50233),
    .O(net_50265)
  );
  InMux inmux_12_11_50235_50279 (
    .I(net_50235),
    .O(net_50279)
  );
  ClkMux inmux_12_11_5_50300 (
    .I(net_5),
    .O(net_50300)
  );
  CEMux inmux_12_12_50345_50422 (
    .I(net_50345),
    .O(net_50422)
  );
  InMux inmux_12_12_50353_50396 (
    .I(net_50353),
    .O(net_50396)
  );
  InMux inmux_12_12_50355_50379 (
    .I(net_50355),
    .O(net_50379)
  );
  InMux inmux_12_12_50362_50394 (
    .I(net_50362),
    .O(net_50394)
  );
  InMux inmux_12_12_50363_50383 (
    .I(net_50363),
    .O(net_50383)
  );
  InMux inmux_12_12_50368_50395 (
    .I(net_50368),
    .O(net_50395)
  );
  InMux inmux_12_12_50372_50397 (
    .I(net_50372),
    .O(net_50397)
  );
  ClkMux inmux_12_12_5_50423 (
    .I(net_5),
    .O(net_50423)
  );
  InMux inmux_12_13_50466_50523 (
    .I(net_50466),
    .O(net_50523)
  );
  InMux inmux_12_13_50472_50532 (
    .I(net_50472),
    .O(net_50532)
  );
  InMux inmux_12_13_50475_50518 (
    .I(net_50475),
    .O(net_50518)
  );
  InMux inmux_12_13_50476_50517 (
    .I(net_50476),
    .O(net_50517)
  );
  InMux inmux_12_13_50477_50501 (
    .I(net_50477),
    .O(net_50501)
  );
  InMux inmux_12_13_50492_50514 (
    .I(net_50492),
    .O(net_50514)
  );
  InMux inmux_12_13_50494_50538 (
    .I(net_50494),
    .O(net_50538)
  );
  ClkMux inmux_12_13_5_50546 (
    .I(net_5),
    .O(net_50546)
  );
  SRMux inmux_12_13_9_50547 (
    .I(net_9),
    .O(net_50547)
  );
  InMux inmux_12_14_50590_50654 (
    .I(net_50590),
    .O(net_50654)
  );
  InMux inmux_12_14_50598_50648 (
    .I(net_50598),
    .O(net_50648)
  );
  InMux inmux_12_14_50599_50649 (
    .I(net_50599),
    .O(net_50649)
  );
  InMux inmux_12_14_50600_50624 (
    .I(net_50600),
    .O(net_50624)
  );
  InMux inmux_12_14_50602_50658 (
    .I(net_50602),
    .O(net_50658)
  );
  InMux inmux_12_14_50606_50625 (
    .I(net_50606),
    .O(net_50625)
  );
  InMux inmux_12_14_50606_50628 (
    .I(net_50606),
    .O(net_50628)
  );
  InMux inmux_12_14_50606_50642 (
    .I(net_50606),
    .O(net_50642)
  );
  InMux inmux_12_14_50606_50647 (
    .I(net_50606),
    .O(net_50647)
  );
  InMux inmux_12_14_50606_50652 (
    .I(net_50606),
    .O(net_50652)
  );
  InMux inmux_12_14_50606_50659 (
    .I(net_50606),
    .O(net_50659)
  );
  InMux inmux_12_14_50609_50643 (
    .I(net_50609),
    .O(net_50643)
  );
  InMux inmux_12_14_50612_50630 (
    .I(net_50612),
    .O(net_50630)
  );
  InMux inmux_12_14_50614_50622 (
    .I(net_50614),
    .O(net_50622)
  );
  InMux inmux_12_14_50616_50629 (
    .I(net_50616),
    .O(net_50629)
  );
  InMux inmux_12_14_50617_50640 (
    .I(net_50617),
    .O(net_50640)
  );
  InMux inmux_12_14_50619_50661 (
    .I(net_50619),
    .O(net_50661)
  );
  ClkMux inmux_12_14_5_50669 (
    .I(net_5),
    .O(net_50669)
  );
  CEMux inmux_12_14_6_50668 (
    .I(net_6),
    .O(net_50668)
  );
  SRMux inmux_12_14_9_50670 (
    .I(net_9),
    .O(net_50670)
  );
  CEMux inmux_12_15_50714_50791 (
    .I(net_50714),
    .O(net_50791)
  );
  InMux inmux_12_15_50715_50765 (
    .I(net_50715),
    .O(net_50765)
  );
  InMux inmux_12_15_50715_50772 (
    .I(net_50715),
    .O(net_50772)
  );
  InMux inmux_12_15_50715_50775 (
    .I(net_50715),
    .O(net_50775)
  );
  InMux inmux_12_15_50715_50787 (
    .I(net_50715),
    .O(net_50787)
  );
  InMux inmux_12_15_50723_50752 (
    .I(net_50723),
    .O(net_50752)
  );
  InMux inmux_12_15_50723_50757 (
    .I(net_50723),
    .O(net_50757)
  );
  InMux inmux_12_15_50724_50748 (
    .I(net_50724),
    .O(net_50748)
  );
  InMux inmux_12_15_50731_50770 (
    .I(net_50731),
    .O(net_50770)
  );
  InMux inmux_12_15_50731_50777 (
    .I(net_50731),
    .O(net_50777)
  );
  InMux inmux_12_15_50734_50766 (
    .I(net_50734),
    .O(net_50766)
  );
  InMux inmux_12_15_50734_50788 (
    .I(net_50734),
    .O(net_50788)
  );
  InMux inmux_12_15_50739_50754 (
    .I(net_50739),
    .O(net_50754)
  );
  InMux inmux_12_15_50739_50759 (
    .I(net_50739),
    .O(net_50759)
  );
  InMux inmux_12_15_50739_50764 (
    .I(net_50739),
    .O(net_50764)
  );
  InMux inmux_12_15_50739_50771 (
    .I(net_50739),
    .O(net_50771)
  );
  InMux inmux_12_15_50739_50776 (
    .I(net_50739),
    .O(net_50776)
  );
  InMux inmux_12_15_50739_50790 (
    .I(net_50739),
    .O(net_50790)
  );
  InMux inmux_12_15_50740_50751 (
    .I(net_50740),
    .O(net_50751)
  );
  InMux inmux_12_15_50740_50760 (
    .I(net_50740),
    .O(net_50760)
  );
  InMux inmux_12_15_50740_50763 (
    .I(net_50740),
    .O(net_50763)
  );
  InMux inmux_12_15_50740_50789 (
    .I(net_50740),
    .O(net_50789)
  );
  InMux inmux_12_15_50742_50753 (
    .I(net_50742),
    .O(net_50753)
  );
  InMux inmux_12_15_50742_50758 (
    .I(net_50742),
    .O(net_50758)
  );
  ClkMux inmux_12_15_5_50792 (
    .I(net_5),
    .O(net_50792)
  );
  SRMux inmux_12_15_9_50793 (
    .I(net_9),
    .O(net_50793)
  );
  InMux inmux_12_16_50835_50880 (
    .I(net_50835),
    .O(net_50880)
  );
  InMux inmux_12_16_50836_50869 (
    .I(net_50836),
    .O(net_50869)
  );
  InMux inmux_12_16_50836_50905 (
    .I(net_50836),
    .O(net_50905)
  );
  InMux inmux_12_16_50837_50901 (
    .I(net_50837),
    .O(net_50901)
  );
  InMux inmux_12_16_50837_50906 (
    .I(net_50837),
    .O(net_50906)
  );
  InMux inmux_12_16_50838_50874 (
    .I(net_50838),
    .O(net_50874)
  );
  InMux inmux_12_16_50838_50910 (
    .I(net_50838),
    .O(net_50910)
  );
  InMux inmux_12_16_50839_50882 (
    .I(net_50839),
    .O(net_50882)
  );
  InMux inmux_12_16_50840_50912 (
    .I(net_50840),
    .O(net_50912)
  );
  InMux inmux_12_16_50841_50877 (
    .I(net_50841),
    .O(net_50877)
  );
  InMux inmux_12_16_50842_50888 (
    .I(net_50842),
    .O(net_50888)
  );
  InMux inmux_12_16_50844_50904 (
    .I(net_50844),
    .O(net_50904)
  );
  InMux inmux_12_16_50846_50868 (
    .I(net_50846),
    .O(net_50868)
  );
  InMux inmux_12_16_50846_50875 (
    .I(net_50846),
    .O(net_50875)
  );
  InMux inmux_12_16_50846_50889 (
    .I(net_50846),
    .O(net_50889)
  );
  InMux inmux_12_16_50846_50899 (
    .I(net_50846),
    .O(net_50899)
  );
  InMux inmux_12_16_50847_50898 (
    .I(net_50847),
    .O(net_50898)
  );
  InMux inmux_12_16_50848_50894 (
    .I(net_50848),
    .O(net_50894)
  );
  InMux inmux_12_16_50849_50871 (
    .I(net_50849),
    .O(net_50871)
  );
  InMux inmux_12_16_50849_50876 (
    .I(net_50849),
    .O(net_50876)
  );
  InMux inmux_12_16_50849_50900 (
    .I(net_50849),
    .O(net_50900)
  );
  InMux inmux_12_16_50850_50870 (
    .I(net_50850),
    .O(net_50870)
  );
  InMux inmux_12_16_50856_50886 (
    .I(net_50856),
    .O(net_50886)
  );
  InMux inmux_12_16_50857_50911 (
    .I(net_50857),
    .O(net_50911)
  );
  InMux inmux_12_16_50858_50907 (
    .I(net_50858),
    .O(net_50907)
  );
  InMux inmux_12_16_50864_50887 (
    .I(net_50864),
    .O(net_50887)
  );
  InMux inmux_12_16_50866_50913 (
    .I(net_50866),
    .O(net_50913)
  );
  ClkMux inmux_12_16_5_50915 (
    .I(net_5),
    .O(net_50915)
  );
  SRMux inmux_12_16_9_50916 (
    .I(net_9),
    .O(net_50916)
  );
  InMux inmux_12_17_50959_51011 (
    .I(net_50959),
    .O(net_51011)
  );
  InMux inmux_12_17_50959_51016 (
    .I(net_50959),
    .O(net_51016)
  );
  InMux inmux_12_17_50966_50999 (
    .I(net_50966),
    .O(net_50999)
  );
  InMux inmux_12_17_50966_51035 (
    .I(net_50966),
    .O(net_51035)
  );
  InMux inmux_12_17_50971_51003 (
    .I(net_50971),
    .O(net_51003)
  );
  InMux inmux_12_17_50978_50993 (
    .I(net_50978),
    .O(net_50993)
  );
  InMux inmux_12_17_50978_51000 (
    .I(net_50978),
    .O(net_51000)
  );
  InMux inmux_12_17_50978_51027 (
    .I(net_50978),
    .O(net_51027)
  );
  InMux inmux_12_17_50996_51006 (
    .I(net_50996),
    .O(net_51006)
  );
  ClkMux inmux_12_17_5_51038 (
    .I(net_5),
    .O(net_51038)
  );
  SRMux inmux_12_17_9_51039 (
    .I(net_9),
    .O(net_51039)
  );
  InMux inmux_12_18_51082_51139 (
    .I(net_51082),
    .O(net_51139)
  );
  CEMux inmux_12_18_51092_51160 (
    .I(net_51092),
    .O(net_51160)
  );
  InMux inmux_12_18_51093_51129 (
    .I(net_51093),
    .O(net_51129)
  );
  ClkMux inmux_12_18_5_51161 (
    .I(net_5),
    .O(net_51161)
  );
  InMux inmux_12_19_51218_51255 (
    .I(net_51218),
    .O(net_51255)
  );
  CEMux inmux_12_19_51231_51283 (
    .I(net_51231),
    .O(net_51283)
  );
  ClkMux inmux_12_19_5_51284 (
    .I(net_5),
    .O(net_51284)
  );
  InMux inmux_12_1_48952_48997 (
    .I(net_48952),
    .O(net_48997)
  );
  InMux inmux_12_1_48954_49009 (
    .I(net_48954),
    .O(net_49009)
  );
  InMux inmux_12_1_48959_48990 (
    .I(net_48959),
    .O(net_48990)
  );
  InMux inmux_12_1_48967_48989 (
    .I(net_48967),
    .O(net_48989)
  );
  InMux inmux_12_1_48967_49001 (
    .I(net_48967),
    .O(net_49001)
  );
  InMux inmux_12_1_48967_49008 (
    .I(net_48967),
    .O(net_49008)
  );
  CEMux inmux_12_1_48968_49029 (
    .I(net_48968),
    .O(net_49029)
  );
  InMux inmux_12_1_48975_48995 (
    .I(net_48975),
    .O(net_48995)
  );
  InMux inmux_12_1_48977_49002 (
    .I(net_48977),
    .O(net_49002)
  );
  InMux inmux_12_1_48979_48985 (
    .I(net_48979),
    .O(net_48985)
  );
  InMux inmux_12_1_48979_48992 (
    .I(net_48979),
    .O(net_48992)
  );
  InMux inmux_12_1_48988_48998 (
    .I(net_48988),
    .O(net_48998)
  );
  InMux inmux_12_1_48994_49004 (
    .I(net_48994),
    .O(net_49004)
  );
  InMux inmux_12_1_49000_49010 (
    .I(net_49000),
    .O(net_49010)
  );
  ClkMux inmux_12_1_5_49030 (
    .I(net_5),
    .O(net_49030)
  );
  SRMux inmux_12_1_9_49031 (
    .I(net_9),
    .O(net_49031)
  );
  InMux inmux_12_2_49115_49148 (
    .I(net_49115),
    .O(net_49148)
  );
  InMux inmux_12_2_49119_49155 (
    .I(net_49119),
    .O(net_49155)
  );
  InMux inmux_12_2_49123_49164 (
    .I(net_49123),
    .O(net_49164)
  );
  InMux inmux_12_2_49124_49158 (
    .I(net_49124),
    .O(net_49158)
  );
  InMux inmux_12_2_49131_49170 (
    .I(net_49131),
    .O(net_49170)
  );
  InMux inmux_12_2_49134_49183 (
    .I(net_49134),
    .O(net_49183)
  );
  ClkMux inmux_12_2_5_49193 (
    .I(net_5),
    .O(net_49193)
  );
  SRMux inmux_12_2_9_49194 (
    .I(net_9),
    .O(net_49194)
  );
  InMux inmux_12_3_49236_49276 (
    .I(net_49236),
    .O(net_49276)
  );
  InMux inmux_12_3_49238_49295 (
    .I(net_49238),
    .O(net_49295)
  );
  InMux inmux_12_3_49239_49289 (
    .I(net_49239),
    .O(net_49289)
  );
  InMux inmux_12_3_49240_49312 (
    .I(net_49240),
    .O(net_49312)
  );
  InMux inmux_12_3_49241_49308 (
    .I(net_49241),
    .O(net_49308)
  );
  InMux inmux_12_3_49246_49282 (
    .I(net_49246),
    .O(net_49282)
  );
  InMux inmux_12_3_49256_49271 (
    .I(net_49256),
    .O(net_49271)
  );
  InMux inmux_12_3_49257_49299 (
    .I(net_49257),
    .O(net_49299)
  );
  InMux inmux_12_3_49258_49314 (
    .I(net_49258),
    .O(net_49314)
  );
  InMux inmux_12_3_49266_49294 (
    .I(net_49266),
    .O(net_49294)
  );
  InMux inmux_12_3_49286_49296 (
    .I(net_49286),
    .O(net_49296)
  );
  ClkMux inmux_12_3_5_49316 (
    .I(net_5),
    .O(net_49316)
  );
  SRMux inmux_12_3_9_49317 (
    .I(net_9),
    .O(net_49317)
  );
  InMux inmux_12_4_49363_49437 (
    .I(net_49363),
    .O(net_49437)
  );
  InMux inmux_12_4_49365_49418 (
    .I(net_49365),
    .O(net_49418)
  );
  InMux inmux_12_4_49366_49405 (
    .I(net_49366),
    .O(net_49405)
  );
  InMux inmux_12_4_49367_49400 (
    .I(net_49367),
    .O(net_49400)
  );
  InMux inmux_12_4_49371_49410 (
    .I(net_49371),
    .O(net_49410)
  );
  InMux inmux_12_4_49373_49398 (
    .I(net_49373),
    .O(net_49398)
  );
  InMux inmux_12_4_49375_49435 (
    .I(net_49375),
    .O(net_49435)
  );
  InMux inmux_12_4_49378_49422 (
    .I(net_49378),
    .O(net_49422)
  );
  InMux inmux_12_4_49379_49428 (
    .I(net_49379),
    .O(net_49428)
  );
  InMux inmux_12_4_49380_49429 (
    .I(net_49380),
    .O(net_49429)
  );
  InMux inmux_12_4_49383_49395 (
    .I(net_49383),
    .O(net_49395)
  );
  InMux inmux_12_4_49384_49399 (
    .I(net_49384),
    .O(net_49399)
  );
  InMux inmux_12_4_49384_49430 (
    .I(net_49384),
    .O(net_49430)
  );
  InMux inmux_12_4_49385_49431 (
    .I(net_49385),
    .O(net_49431)
  );
  CEMux inmux_12_4_49386_49438 (
    .I(net_49386),
    .O(net_49438)
  );
  InMux inmux_12_4_49388_49401 (
    .I(net_49388),
    .O(net_49401)
  );
  InMux inmux_12_4_49390_49425 (
    .I(net_49390),
    .O(net_49425)
  );
  ClkMux inmux_12_4_5_49439 (
    .I(net_5),
    .O(net_49439)
  );
  CEMux inmux_12_5_12_49561 (
    .I(net_12),
    .O(net_49561)
  );
  InMux inmux_12_5_49493_49527 (
    .I(net_49493),
    .O(net_49527)
  );
  InMux inmux_12_5_49494_49552 (
    .I(net_49494),
    .O(net_49552)
  );
  InMux inmux_12_5_49495_49517 (
    .I(net_49495),
    .O(net_49517)
  );
  InMux inmux_12_5_49511_49546 (
    .I(net_49511),
    .O(net_49546)
  );
  ClkMux inmux_12_5_5_49562 (
    .I(net_5),
    .O(net_49562)
  );
  InMux inmux_12_6_49608_49665 (
    .I(net_49608),
    .O(net_49665)
  );
  InMux inmux_12_6_49610_49663 (
    .I(net_49610),
    .O(net_49663)
  );
  InMux inmux_12_6_49610_49670 (
    .I(net_49610),
    .O(net_49670)
  );
  InMux inmux_12_6_49610_49677 (
    .I(net_49610),
    .O(net_49677)
  );
  InMux inmux_12_6_49616_49683 (
    .I(net_49616),
    .O(net_49683)
  );
  InMux inmux_12_6_49617_49656 (
    .I(net_49617),
    .O(net_49656)
  );
  InMux inmux_12_6_49620_49640 (
    .I(net_49620),
    .O(net_49640)
  );
  InMux inmux_12_6_49623_49645 (
    .I(net_49623),
    .O(net_49645)
  );
  InMux inmux_12_6_49629_49653 (
    .I(net_49629),
    .O(net_49653)
  );
  InMux inmux_12_6_49630_49671 (
    .I(net_49630),
    .O(net_49671)
  );
  InMux inmux_12_6_49636_49674 (
    .I(net_49636),
    .O(net_49674)
  );
  ClkMux inmux_12_6_5_49685 (
    .I(net_5),
    .O(net_49685)
  );
  SRMux inmux_12_6_9_49686 (
    .I(net_9),
    .O(net_49686)
  );
  InMux inmux_12_7_49737_49780 (
    .I(net_49737),
    .O(net_49780)
  );
  InMux inmux_12_7_49739_49763 (
    .I(net_49739),
    .O(net_49763)
  );
  InMux inmux_12_7_49741_49785 (
    .I(net_49741),
    .O(net_49785)
  );
  InMux inmux_12_7_49742_49781 (
    .I(net_49742),
    .O(net_49781)
  );
  InMux inmux_12_7_49744_49804 (
    .I(net_49744),
    .O(net_49804)
  );
  InMux inmux_12_7_49745_49779 (
    .I(net_49745),
    .O(net_49779)
  );
  InMux inmux_12_7_49750_49797 (
    .I(net_49750),
    .O(net_49797)
  );
  InMux inmux_12_7_49752_49767 (
    .I(net_49752),
    .O(net_49767)
  );
  InMux inmux_12_7_49755_49782 (
    .I(net_49755),
    .O(net_49782)
  );
  ClkMux inmux_12_7_5_49808 (
    .I(net_5),
    .O(net_49808)
  );
  CEMux inmux_12_7_8_49807 (
    .I(net_8),
    .O(net_49807)
  );
  CEMux inmux_12_8_10_49930 (
    .I(net_10),
    .O(net_49930)
  );
  InMux inmux_12_8_49855_49886 (
    .I(net_49855),
    .O(net_49886)
  );
  InMux inmux_12_8_49857_49927 (
    .I(net_49857),
    .O(net_49927)
  );
  InMux inmux_12_8_49859_49909 (
    .I(net_49859),
    .O(net_49909)
  );
  InMux inmux_12_8_49861_49916 (
    .I(net_49861),
    .O(net_49916)
  );
  ClkMux inmux_12_8_5_49931 (
    .I(net_5),
    .O(net_49931)
  );
  InMux inmux_12_9_49985_50038 (
    .I(net_49985),
    .O(net_50038)
  );
  InMux inmux_12_9_49993_50010 (
    .I(net_49993),
    .O(net_50010)
  );
  InMux inmux_12_9_49998_50046 (
    .I(net_49998),
    .O(net_50046)
  );
  CEMux inmux_12_9_50001_50053 (
    .I(net_50001),
    .O(net_50053)
  );
  ClkMux inmux_12_9_5_50054 (
    .I(net_5),
    .O(net_50054)
  );
  InMux inmux_13_10_53929_53974 (
    .I(net_53929),
    .O(net_53974)
  );
  InMux inmux_13_10_53940_53962 (
    .I(net_53940),
    .O(net_53962)
  );
  InMux inmux_13_10_53940_53988 (
    .I(net_53940),
    .O(net_53988)
  );
  InMux inmux_13_10_53941_53987 (
    .I(net_53941),
    .O(net_53987)
  );
  InMux inmux_13_10_53942_53964 (
    .I(net_53942),
    .O(net_53964)
  );
  InMux inmux_13_10_53944_53961 (
    .I(net_53944),
    .O(net_53961)
  );
  InMux inmux_13_10_53945_53969 (
    .I(net_53945),
    .O(net_53969)
  );
  InMux inmux_13_10_53946_53985 (
    .I(net_53946),
    .O(net_53985)
  );
  InMux inmux_13_10_53949_53991 (
    .I(net_53949),
    .O(net_53991)
  );
  InMux inmux_13_10_53952_53986 (
    .I(net_53952),
    .O(net_53986)
  );
  InMux inmux_13_10_53953_53963 (
    .I(net_53953),
    .O(net_53963)
  );
  CEMux inmux_13_10_53955_54007 (
    .I(net_53955),
    .O(net_54007)
  );
  ClkMux inmux_13_10_5_54008 (
    .I(net_5),
    .O(net_54008)
  );
  InMux inmux_13_11_54055_54108 (
    .I(net_54055),
    .O(net_54108)
  );
  InMux inmux_13_11_54056_54109 (
    .I(net_54056),
    .O(net_54109)
  );
  InMux inmux_13_11_54058_54116 (
    .I(net_54058),
    .O(net_54116)
  );
  InMux inmux_13_11_54066_54093 (
    .I(net_54066),
    .O(net_54093)
  );
  InMux inmux_13_11_54070_54099 (
    .I(net_54070),
    .O(net_54099)
  );
  InMux inmux_13_11_54072_54111 (
    .I(net_54072),
    .O(net_54111)
  );
  InMux inmux_13_11_54073_54110 (
    .I(net_54073),
    .O(net_54110)
  );
  CEMux inmux_13_11_54078_54130 (
    .I(net_54078),
    .O(net_54130)
  );
  InMux inmux_13_11_54082_54122 (
    .I(net_54082),
    .O(net_54122)
  );
  ClkMux inmux_13_11_5_54131 (
    .I(net_5),
    .O(net_54131)
  );
  CEMux inmux_13_12_54176_54253 (
    .I(net_54176),
    .O(net_54253)
  );
  InMux inmux_13_12_54179_54220 (
    .I(net_54179),
    .O(net_54220)
  );
  InMux inmux_13_12_54180_54216 (
    .I(net_54180),
    .O(net_54216)
  );
  InMux inmux_13_12_54183_54245 (
    .I(net_54183),
    .O(net_54245)
  );
  InMux inmux_13_12_54184_54251 (
    .I(net_54184),
    .O(net_54251)
  );
  InMux inmux_13_12_54195_54232 (
    .I(net_54195),
    .O(net_54232)
  );
  InMux inmux_13_12_54196_54207 (
    .I(net_54196),
    .O(net_54207)
  );
  InMux inmux_13_12_54199_54228 (
    .I(net_54199),
    .O(net_54228)
  );
  InMux inmux_13_12_54205_54240 (
    .I(net_54205),
    .O(net_54240)
  );
  ClkMux inmux_13_12_5_54254 (
    .I(net_5),
    .O(net_54254)
  );
  InMux inmux_13_13_54299_54337 (
    .I(net_54299),
    .O(net_54337)
  );
  InMux inmux_13_13_54299_54354 (
    .I(net_54299),
    .O(net_54354)
  );
  InMux inmux_13_13_54299_54366 (
    .I(net_54299),
    .O(net_54366)
  );
  InMux inmux_13_13_54299_54375 (
    .I(net_54299),
    .O(net_54375)
  );
  InMux inmux_13_13_54303_54373 (
    .I(net_54303),
    .O(net_54373)
  );
  InMux inmux_13_13_54304_54360 (
    .I(net_54304),
    .O(net_54360)
  );
  InMux inmux_13_13_54305_54355 (
    .I(net_54305),
    .O(net_54355)
  );
  InMux inmux_13_13_54307_54369 (
    .I(net_54307),
    .O(net_54369)
  );
  InMux inmux_13_13_54308_54339 (
    .I(net_54308),
    .O(net_54339)
  );
  InMux inmux_13_13_54309_54345 (
    .I(net_54309),
    .O(net_54345)
  );
  InMux inmux_13_13_54311_54336 (
    .I(net_54311),
    .O(net_54336)
  );
  InMux inmux_13_13_54311_54357 (
    .I(net_54311),
    .O(net_54357)
  );
  InMux inmux_13_13_54311_54367 (
    .I(net_54311),
    .O(net_54367)
  );
  InMux inmux_13_13_54311_54374 (
    .I(net_54311),
    .O(net_54374)
  );
  InMux inmux_13_13_54313_54356 (
    .I(net_54313),
    .O(net_54356)
  );
  InMux inmux_13_13_54316_54372 (
    .I(net_54316),
    .O(net_54372)
  );
  InMux inmux_13_13_54317_54351 (
    .I(net_54317),
    .O(net_54351)
  );
  InMux inmux_13_13_54323_54338 (
    .I(net_54323),
    .O(net_54338)
  );
  CEMux inmux_13_13_54324_54376 (
    .I(net_54324),
    .O(net_54376)
  );
  InMux inmux_13_13_54325_54331 (
    .I(net_54325),
    .O(net_54331)
  );
  InMux inmux_13_13_54326_54368 (
    .I(net_54326),
    .O(net_54368)
  );
  ClkMux inmux_13_13_5_54377 (
    .I(net_5),
    .O(net_54377)
  );
  InMux inmux_13_14_54425_54478 (
    .I(net_54425),
    .O(net_54478)
  );
  InMux inmux_13_14_54427_54461 (
    .I(net_54427),
    .O(net_54461)
  );
  InMux inmux_13_14_54428_54495 (
    .I(net_54428),
    .O(net_54495)
  );
  InMux inmux_13_14_54429_54453 (
    .I(net_54429),
    .O(net_54453)
  );
  InMux inmux_13_14_54431_54496 (
    .I(net_54431),
    .O(net_54496)
  );
  InMux inmux_13_14_54433_54491 (
    .I(net_54433),
    .O(net_54491)
  );
  InMux inmux_13_14_54435_54498 (
    .I(net_54435),
    .O(net_54498)
  );
  InMux inmux_13_14_54436_54486 (
    .I(net_54436),
    .O(net_54486)
  );
  InMux inmux_13_14_54437_54471 (
    .I(net_54437),
    .O(net_54471)
  );
  InMux inmux_13_14_54438_54465 (
    .I(net_54438),
    .O(net_54465)
  );
  InMux inmux_13_14_54444_54459 (
    .I(net_54444),
    .O(net_54459)
  );
  InMux inmux_13_14_54446_54497 (
    .I(net_54446),
    .O(net_54497)
  );
  CEMux inmux_13_14_54447_54499 (
    .I(net_54447),
    .O(net_54499)
  );
  InMux inmux_13_14_54450_54466 (
    .I(net_54450),
    .O(net_54466)
  );
  ClkMux inmux_13_14_5_54500 (
    .I(net_5),
    .O(net_54500)
  );
  InMux inmux_13_15_54543_54607 (
    .I(net_54543),
    .O(net_54607)
  );
  InMux inmux_13_15_54544_54584 (
    .I(net_54544),
    .O(net_54584)
  );
  InMux inmux_13_15_54544_54589 (
    .I(net_54544),
    .O(net_54589)
  );
  InMux inmux_13_15_54546_54582 (
    .I(net_54546),
    .O(net_54582)
  );
  InMux inmux_13_15_54549_54588 (
    .I(net_54549),
    .O(net_54588)
  );
  InMux inmux_13_15_54551_54615 (
    .I(net_54551),
    .O(net_54615)
  );
  InMux inmux_13_15_54552_54578 (
    .I(net_54552),
    .O(net_54578)
  );
  InMux inmux_13_15_54553_54620 (
    .I(net_54553),
    .O(net_54620)
  );
  CEMux inmux_13_15_54554_54622 (
    .I(net_54554),
    .O(net_54622)
  );
  InMux inmux_13_15_54555_54591 (
    .I(net_54555),
    .O(net_54591)
  );
  InMux inmux_13_15_54556_54585 (
    .I(net_54556),
    .O(net_54585)
  );
  InMux inmux_13_15_54561_54576 (
    .I(net_54561),
    .O(net_54576)
  );
  InMux inmux_13_15_54567_54603 (
    .I(net_54567),
    .O(net_54603)
  );
  InMux inmux_13_15_54574_54590 (
    .I(net_54574),
    .O(net_54590)
  );
  ClkMux inmux_13_15_5_54623 (
    .I(net_5),
    .O(net_54623)
  );
  InMux inmux_13_16_54667_54707 (
    .I(net_54667),
    .O(net_54707)
  );
  InMux inmux_13_16_54668_54730 (
    .I(net_54668),
    .O(net_54730)
  );
  InMux inmux_13_16_54668_54737 (
    .I(net_54668),
    .O(net_54737)
  );
  InMux inmux_13_16_54669_54700 (
    .I(net_54669),
    .O(net_54700)
  );
  InMux inmux_13_16_54670_54735 (
    .I(net_54670),
    .O(net_54735)
  );
  InMux inmux_13_16_54672_54723 (
    .I(net_54672),
    .O(net_54723)
  );
  InMux inmux_13_16_54673_54729 (
    .I(net_54673),
    .O(net_54729)
  );
  InMux inmux_13_16_54676_54726 (
    .I(net_54676),
    .O(net_54726)
  );
  InMux inmux_13_16_54677_54708 (
    .I(net_54677),
    .O(net_54708)
  );
  InMux inmux_13_16_54678_54738 (
    .I(net_54678),
    .O(net_54738)
  );
  InMux inmux_13_16_54679_54725 (
    .I(net_54679),
    .O(net_54725)
  );
  InMux inmux_13_16_54682_54720 (
    .I(net_54682),
    .O(net_54720)
  );
  InMux inmux_13_16_54685_54731 (
    .I(net_54685),
    .O(net_54731)
  );
  InMux inmux_13_16_54694_54719 (
    .I(net_54694),
    .O(net_54719)
  );
  InMux inmux_13_16_54694_54724 (
    .I(net_54694),
    .O(net_54724)
  );
  InMux inmux_13_16_54695_54711 (
    .I(net_54695),
    .O(net_54711)
  );
  InMux inmux_13_16_54695_54742 (
    .I(net_54695),
    .O(net_54742)
  );
  InMux inmux_13_16_54696_54736 (
    .I(net_54696),
    .O(net_54736)
  );
  InMux inmux_13_16_54704_54714 (
    .I(net_54704),
    .O(net_54714)
  );
  ClkMux inmux_13_16_5_54746 (
    .I(net_5),
    .O(net_54746)
  );
  SRMux inmux_13_16_9_54747 (
    .I(net_9),
    .O(net_54747)
  );
  InMux inmux_13_17_54789_54853 (
    .I(net_54789),
    .O(net_54853)
  );
  InMux inmux_13_17_54790_54842 (
    .I(net_54790),
    .O(net_54842)
  );
  InMux inmux_13_17_54790_54847 (
    .I(net_54790),
    .O(net_54847)
  );
  InMux inmux_13_17_54793_54831 (
    .I(net_54793),
    .O(net_54831)
  );
  InMux inmux_13_17_54796_54828 (
    .I(net_54796),
    .O(net_54828)
  );
  InMux inmux_13_17_54796_54854 (
    .I(net_54796),
    .O(net_54854)
  );
  InMux inmux_13_17_54800_54829 (
    .I(net_54800),
    .O(net_54829)
  );
  InMux inmux_13_17_54803_54852 (
    .I(net_54803),
    .O(net_54852)
  );
  InMux inmux_13_17_54804_54855 (
    .I(net_54804),
    .O(net_54855)
  );
  InMux inmux_13_17_54816_54865 (
    .I(net_54816),
    .O(net_54865)
  );
  ClkMux inmux_13_17_5_54869 (
    .I(net_5),
    .O(net_54869)
  );
  SRMux inmux_13_17_9_54870 (
    .I(net_9),
    .O(net_54870)
  );
  InMux inmux_13_18_54912_54959 (
    .I(net_54912),
    .O(net_54959)
  );
  InMux inmux_13_18_54913_54946 (
    .I(net_54913),
    .O(net_54946)
  );
  InMux inmux_13_18_54915_54958 (
    .I(net_54915),
    .O(net_54958)
  );
  InMux inmux_13_18_54916_54978 (
    .I(net_54916),
    .O(net_54978)
  );
  InMux inmux_13_18_54917_54989 (
    .I(net_54917),
    .O(net_54989)
  );
  InMux inmux_13_18_54919_54987 (
    .I(net_54919),
    .O(net_54987)
  );
  InMux inmux_13_18_54920_54963 (
    .I(net_54920),
    .O(net_54963)
  );
  CEMux inmux_13_18_54923_54991 (
    .I(net_54923),
    .O(net_54991)
  );
  InMux inmux_13_18_54924_54953 (
    .I(net_54924),
    .O(net_54953)
  );
  InMux inmux_13_18_54925_54981 (
    .I(net_54925),
    .O(net_54981)
  );
  InMux inmux_13_18_54926_54984 (
    .I(net_54926),
    .O(net_54984)
  );
  InMux inmux_13_18_54927_54947 (
    .I(net_54927),
    .O(net_54947)
  );
  InMux inmux_13_18_54927_54954 (
    .I(net_54927),
    .O(net_54954)
  );
  InMux inmux_13_18_54927_54957 (
    .I(net_54927),
    .O(net_54957)
  );
  InMux inmux_13_18_54927_54964 (
    .I(net_54927),
    .O(net_54964)
  );
  InMux inmux_13_18_54927_54976 (
    .I(net_54927),
    .O(net_54976)
  );
  InMux inmux_13_18_54927_54983 (
    .I(net_54927),
    .O(net_54983)
  );
  InMux inmux_13_18_54927_54988 (
    .I(net_54927),
    .O(net_54988)
  );
  InMux inmux_13_18_54928_54966 (
    .I(net_54928),
    .O(net_54966)
  );
  InMux inmux_13_18_54929_54951 (
    .I(net_54929),
    .O(net_54951)
  );
  InMux inmux_13_18_54930_54952 (
    .I(net_54930),
    .O(net_54952)
  );
  InMux inmux_13_18_54931_54960 (
    .I(net_54931),
    .O(net_54960)
  );
  InMux inmux_13_18_54933_54975 (
    .I(net_54933),
    .O(net_54975)
  );
  InMux inmux_13_18_54935_54948 (
    .I(net_54935),
    .O(net_54948)
  );
  InMux inmux_13_18_54936_54977 (
    .I(net_54936),
    .O(net_54977)
  );
  InMux inmux_13_18_54938_54965 (
    .I(net_54938),
    .O(net_54965)
  );
  InMux inmux_13_18_54939_54945 (
    .I(net_54939),
    .O(net_54945)
  );
  InMux inmux_13_18_54941_54990 (
    .I(net_54941),
    .O(net_54990)
  );
  InMux inmux_13_18_54942_54982 (
    .I(net_54942),
    .O(net_54982)
  );
  ClkMux inmux_13_18_5_54992 (
    .I(net_5),
    .O(net_54992)
  );
  InMux inmux_13_19_55036_55110 (
    .I(net_55036),
    .O(net_55110)
  );
  InMux inmux_13_19_55039_55113 (
    .I(net_55039),
    .O(net_55113)
  );
  InMux inmux_13_19_55044_55111 (
    .I(net_55044),
    .O(net_55111)
  );
  CEMux inmux_13_19_55046_55114 (
    .I(net_55046),
    .O(net_55114)
  );
  InMux inmux_13_19_55049_55112 (
    .I(net_55049),
    .O(net_55112)
  );
  ClkMux inmux_13_19_5_55115 (
    .I(net_5),
    .O(net_55115)
  );
  InMux inmux_13_1_52784_52846 (
    .I(net_52784),
    .O(net_52846)
  );
  InMux inmux_13_1_52785_52850 (
    .I(net_52785),
    .O(net_52850)
  );
  InMux inmux_13_1_52791_52851 (
    .I(net_52791),
    .O(net_52851)
  );
  InMux inmux_13_1_52792_52847 (
    .I(net_52792),
    .O(net_52847)
  );
  InMux inmux_13_1_52792_52852 (
    .I(net_52792),
    .O(net_52852)
  );
  InMux inmux_13_1_52793_52832 (
    .I(net_52793),
    .O(net_52832)
  );
  ClkMux inmux_13_1_5_52861 (
    .I(net_5),
    .O(net_52861)
  );
  SRMux inmux_13_1_9_52862 (
    .I(net_9),
    .O(net_52862)
  );
  InMux inmux_13_2_52948_52977 (
    .I(net_52948),
    .O(net_52977)
  );
  InMux inmux_13_2_52948_52998 (
    .I(net_52948),
    .O(net_52998)
  );
  InMux inmux_13_2_52952_53002 (
    .I(net_52952),
    .O(net_53002)
  );
  InMux inmux_13_2_52954_52980 (
    .I(net_52954),
    .O(net_52980)
  );
  InMux inmux_13_2_52954_52995 (
    .I(net_52954),
    .O(net_52995)
  );
  CEMux inmux_13_2_52955_53023 (
    .I(net_52955),
    .O(net_53023)
  );
  InMux inmux_13_2_52959_52986 (
    .I(net_52959),
    .O(net_52986)
  );
  InMux inmux_13_2_52963_52990 (
    .I(net_52963),
    .O(net_52990)
  );
  InMux inmux_13_2_52970_52985 (
    .I(net_52970),
    .O(net_52985)
  );
  InMux inmux_13_2_52971_52984 (
    .I(net_52971),
    .O(net_52984)
  );
  ClkMux inmux_13_2_5_53024 (
    .I(net_5),
    .O(net_53024)
  );
  SRMux inmux_13_2_9_53025 (
    .I(net_9),
    .O(net_53025)
  );
  IoInMux inmux_13_31_56527_56518 (
    .I(net_56527),
    .O(net_56518)
  );
  IoInMux inmux_13_31_56533_56515 (
    .I(net_56533),
    .O(net_56515)
  );
  InMux inmux_13_3_53067_53138 (
    .I(net_53067),
    .O(net_53138)
  );
  InMux inmux_13_3_53068_53142 (
    .I(net_53068),
    .O(net_53142)
  );
  InMux inmux_13_3_53070_53144 (
    .I(net_53070),
    .O(net_53144)
  );
  InMux inmux_13_3_53073_53131 (
    .I(net_53073),
    .O(net_53131)
  );
  InMux inmux_13_3_53074_53101 (
    .I(net_53074),
    .O(net_53101)
  );
  InMux inmux_13_3_53080_53145 (
    .I(net_53080),
    .O(net_53145)
  );
  InMux inmux_13_3_53083_53109 (
    .I(net_53083),
    .O(net_53109)
  );
  InMux inmux_13_3_53087_53112 (
    .I(net_53087),
    .O(net_53112)
  );
  InMux inmux_13_3_53088_53127 (
    .I(net_53088),
    .O(net_53127)
  );
  InMux inmux_13_3_53092_53126 (
    .I(net_53092),
    .O(net_53126)
  );
  InMux inmux_13_3_53093_53132 (
    .I(net_53093),
    .O(net_53132)
  );
  ClkMux inmux_13_3_5_53147 (
    .I(net_5),
    .O(net_53147)
  );
  SRMux inmux_13_3_9_53148 (
    .I(net_9),
    .O(net_53148)
  );
  InMux inmux_13_4_53192_53259 (
    .I(net_53192),
    .O(net_53259)
  );
  InMux inmux_13_4_53193_53262 (
    .I(net_53193),
    .O(net_53262)
  );
  InMux inmux_13_4_53194_53261 (
    .I(net_53194),
    .O(net_53261)
  );
  InMux inmux_13_4_53195_53231 (
    .I(net_53195),
    .O(net_53231)
  );
  InMux inmux_13_4_53198_53260 (
    .I(net_53198),
    .O(net_53260)
  );
  InMux inmux_13_4_53199_53244 (
    .I(net_53199),
    .O(net_53244)
  );
  InMux inmux_13_4_53200_53265 (
    .I(net_53200),
    .O(net_53265)
  );
  InMux inmux_13_4_53201_53242 (
    .I(net_53201),
    .O(net_53242)
  );
  InMux inmux_13_4_53203_53223 (
    .I(net_53203),
    .O(net_53223)
  );
  InMux inmux_13_4_53206_53256 (
    .I(net_53206),
    .O(net_53256)
  );
  InMux inmux_13_4_53207_53248 (
    .I(net_53207),
    .O(net_53248)
  );
  InMux inmux_13_4_53210_53268 (
    .I(net_53210),
    .O(net_53268)
  );
  InMux inmux_13_4_53211_53241 (
    .I(net_53211),
    .O(net_53241)
  );
  InMux inmux_13_4_53217_53235 (
    .I(net_53217),
    .O(net_53235)
  );
  ClkMux inmux_13_4_5_53270 (
    .I(net_5),
    .O(net_53270)
  );
  SRMux inmux_13_4_9_53271 (
    .I(net_9),
    .O(net_53271)
  );
  InMux inmux_13_5_53315_53346 (
    .I(net_53315),
    .O(net_53346)
  );
  InMux inmux_13_5_53322_53377 (
    .I(net_53322),
    .O(net_53377)
  );
  CEMux inmux_13_5_53324_53392 (
    .I(net_53324),
    .O(net_53392)
  );
  InMux inmux_13_5_53331_53384 (
    .I(net_53331),
    .O(net_53384)
  );
  InMux inmux_13_5_53332_53354 (
    .I(net_53332),
    .O(net_53354)
  );
  ClkMux inmux_13_5_5_53393 (
    .I(net_5),
    .O(net_53393)
  );
  CEMux inmux_13_6_12_53515 (
    .I(net_12),
    .O(net_53515)
  );
  InMux inmux_13_6_53439_53484 (
    .I(net_53439),
    .O(net_53484)
  );
  InMux inmux_13_6_53441_53472 (
    .I(net_53441),
    .O(net_53472)
  );
  InMux inmux_13_6_53445_53493 (
    .I(net_53445),
    .O(net_53493)
  );
  InMux inmux_13_6_53450_53487 (
    .I(net_53450),
    .O(net_53487)
  );
  InMux inmux_13_6_53451_53500 (
    .I(net_53451),
    .O(net_53500)
  );
  InMux inmux_13_6_53453_53496 (
    .I(net_53453),
    .O(net_53496)
  );
  InMux inmux_13_6_53454_53505 (
    .I(net_53454),
    .O(net_53505)
  );
  InMux inmux_13_6_53455_53475 (
    .I(net_53455),
    .O(net_53475)
  );
  InMux inmux_13_6_53458_53495 (
    .I(net_53458),
    .O(net_53495)
  );
  InMux inmux_13_6_53462_53494 (
    .I(net_53462),
    .O(net_53494)
  );
  InMux inmux_13_6_53467_53512 (
    .I(net_53467),
    .O(net_53512)
  );
  ClkMux inmux_13_6_5_53516 (
    .I(net_5),
    .O(net_53516)
  );
  InMux inmux_13_7_53559_53606 (
    .I(net_53559),
    .O(net_53606)
  );
  InMux inmux_13_7_53564_53600 (
    .I(net_53564),
    .O(net_53600)
  );
  InMux inmux_13_7_53566_53634 (
    .I(net_53566),
    .O(net_53634)
  );
  InMux inmux_13_7_53567_53595 (
    .I(net_53567),
    .O(net_53595)
  );
  InMux inmux_13_7_53569_53636 (
    .I(net_53569),
    .O(net_53636)
  );
  CEMux inmux_13_7_53570_53638 (
    .I(net_53570),
    .O(net_53638)
  );
  InMux inmux_13_7_53578_53610 (
    .I(net_53578),
    .O(net_53610)
  );
  InMux inmux_13_7_53579_53637 (
    .I(net_53579),
    .O(net_53637)
  );
  InMux inmux_13_7_53580_53605 (
    .I(net_53580),
    .O(net_53605)
  );
  InMux inmux_13_7_53584_53630 (
    .I(net_53584),
    .O(net_53630)
  );
  InMux inmux_13_7_53586_53635 (
    .I(net_53586),
    .O(net_53635)
  );
  InMux inmux_13_7_53587_53607 (
    .I(net_53587),
    .O(net_53607)
  );
  InMux inmux_13_7_53588_53604 (
    .I(net_53588),
    .O(net_53604)
  );
  InMux inmux_13_7_53589_53624 (
    .I(net_53589),
    .O(net_53624)
  );
  InMux inmux_13_7_53590_53616 (
    .I(net_53590),
    .O(net_53616)
  );
  ClkMux inmux_13_7_5_53639 (
    .I(net_5),
    .O(net_53639)
  );
  InMux inmux_13_8_53682_53727 (
    .I(net_53682),
    .O(net_53727)
  );
  InMux inmux_13_8_53682_53741 (
    .I(net_53682),
    .O(net_53741)
  );
  InMux inmux_13_8_53682_53746 (
    .I(net_53682),
    .O(net_53746)
  );
  InMux inmux_13_8_53682_53751 (
    .I(net_53682),
    .O(net_53751)
  );
  InMux inmux_13_8_53682_53758 (
    .I(net_53682),
    .O(net_53758)
  );
  InMux inmux_13_8_53684_53715 (
    .I(net_53684),
    .O(net_53715)
  );
  InMux inmux_13_8_53685_53747 (
    .I(net_53685),
    .O(net_53747)
  );
  InMux inmux_13_8_53686_53739 (
    .I(net_53686),
    .O(net_53739)
  );
  InMux inmux_13_8_53687_53718 (
    .I(net_53687),
    .O(net_53718)
  );
  InMux inmux_13_8_53687_53721 (
    .I(net_53687),
    .O(net_53721)
  );
  InMux inmux_13_8_53688_53717 (
    .I(net_53688),
    .O(net_53717)
  );
  InMux inmux_13_8_53691_53753 (
    .I(net_53691),
    .O(net_53753)
  );
  InMux inmux_13_8_53692_53754 (
    .I(net_53692),
    .O(net_53754)
  );
  InMux inmux_13_8_53693_53724 (
    .I(net_53693),
    .O(net_53724)
  );
  InMux inmux_13_8_53695_53722 (
    .I(net_53695),
    .O(net_53722)
  );
  InMux inmux_13_8_53696_53745 (
    .I(net_53696),
    .O(net_53745)
  );
  InMux inmux_13_8_53699_53728 (
    .I(net_53699),
    .O(net_53728)
  );
  InMux inmux_13_8_53701_53716 (
    .I(net_53701),
    .O(net_53716)
  );
  InMux inmux_13_8_53701_53723 (
    .I(net_53701),
    .O(net_53723)
  );
  InMux inmux_13_8_53702_53760 (
    .I(net_53702),
    .O(net_53760)
  );
  InMux inmux_13_8_53703_53757 (
    .I(net_53703),
    .O(net_53757)
  );
  InMux inmux_13_8_53711_53729 (
    .I(net_53711),
    .O(net_53729)
  );
  InMux inmux_13_8_53712_53742 (
    .I(net_53712),
    .O(net_53742)
  );
  ClkMux inmux_13_8_5_53762 (
    .I(net_5),
    .O(net_53762)
  );
  CEMux inmux_13_8_6_53761 (
    .I(net_6),
    .O(net_53761)
  );
  SRMux inmux_13_8_9_53763 (
    .I(net_9),
    .O(net_53763)
  );
  InMux inmux_13_9_53811_53852 (
    .I(net_53811),
    .O(net_53852)
  );
  InMux inmux_13_9_53816_53871 (
    .I(net_53816),
    .O(net_53871)
  );
  CEMux inmux_13_9_53832_53884 (
    .I(net_53832),
    .O(net_53884)
  );
  ClkMux inmux_13_9_5_53885 (
    .I(net_5),
    .O(net_53885)
  );
  InMux inmux_14_10_57759_57792 (
    .I(net_57759),
    .O(net_57792)
  );
  InMux inmux_14_10_57759_57797 (
    .I(net_57759),
    .O(net_57797)
  );
  InMux inmux_14_10_57759_57804 (
    .I(net_57759),
    .O(net_57804)
  );
  InMux inmux_14_10_57759_57809 (
    .I(net_57759),
    .O(net_57809)
  );
  InMux inmux_14_10_57759_57821 (
    .I(net_57759),
    .O(net_57821)
  );
  InMux inmux_14_10_57759_57828 (
    .I(net_57759),
    .O(net_57828)
  );
  InMux inmux_14_10_57759_57835 (
    .I(net_57759),
    .O(net_57835)
  );
  InMux inmux_14_10_57760_57803 (
    .I(net_57760),
    .O(net_57803)
  );
  InMux inmux_14_10_57771_57834 (
    .I(net_57771),
    .O(net_57834)
  );
  InMux inmux_14_10_57773_57824 (
    .I(net_57773),
    .O(net_57824)
  );
  InMux inmux_14_10_57774_57817 (
    .I(net_57774),
    .O(net_57817)
  );
  InMux inmux_14_10_57778_57810 (
    .I(net_57778),
    .O(net_57810)
  );
  InMux inmux_14_10_57781_57799 (
    .I(net_57781),
    .O(net_57799)
  );
  InMux inmux_14_10_57782_57794 (
    .I(net_57782),
    .O(net_57794)
  );
  InMux inmux_14_10_57786_57830 (
    .I(net_57786),
    .O(net_57830)
  );
  ClkMux inmux_14_10_5_57838 (
    .I(net_5),
    .O(net_57838)
  );
  SRMux inmux_14_10_9_57839 (
    .I(net_9),
    .O(net_57839)
  );
  CEMux inmux_14_11_57883_57960 (
    .I(net_57883),
    .O(net_57960)
  );
  InMux inmux_14_11_57884_57939 (
    .I(net_57884),
    .O(net_57939)
  );
  InMux inmux_14_11_57890_57914 (
    .I(net_57890),
    .O(net_57914)
  );
  InMux inmux_14_11_57893_57934 (
    .I(net_57893),
    .O(net_57934)
  );
  InMux inmux_14_11_57896_57959 (
    .I(net_57896),
    .O(net_57959)
  );
  ClkMux inmux_14_11_5_57961 (
    .I(net_5),
    .O(net_57961)
  );
  InMux inmux_14_12_58012_58062 (
    .I(net_58012),
    .O(net_58062)
  );
  ClkMux inmux_14_12_5_58084 (
    .I(net_5),
    .O(net_58084)
  );
  SRMux inmux_14_12_9_58085 (
    .I(net_9),
    .O(net_58085)
  );
  InMux inmux_14_13_58131_58193 (
    .I(net_58131),
    .O(net_58193)
  );
  InMux inmux_14_13_58133_58198 (
    .I(net_58133),
    .O(net_58198)
  );
  InMux inmux_14_13_58139_58180 (
    .I(net_58139),
    .O(net_58180)
  );
  InMux inmux_14_13_58139_58199 (
    .I(net_58139),
    .O(net_58199)
  );
  InMux inmux_14_13_58143_58167 (
    .I(net_58143),
    .O(net_58167)
  );
  InMux inmux_14_13_58144_58204 (
    .I(net_58144),
    .O(net_58204)
  );
  InMux inmux_14_13_58145_58174 (
    .I(net_58145),
    .O(net_58174)
  );
  InMux inmux_14_13_58147_58186 (
    .I(net_58147),
    .O(net_58186)
  );
  InMux inmux_14_13_58151_58178 (
    .I(net_58151),
    .O(net_58178)
  );
  InMux inmux_14_13_58152_58160 (
    .I(net_58152),
    .O(net_58160)
  );
  InMux inmux_14_13_58154_58179 (
    .I(net_58154),
    .O(net_58179)
  );
  InMux inmux_14_13_58154_58196 (
    .I(net_58154),
    .O(net_58196)
  );
  InMux inmux_14_13_58155_58197 (
    .I(net_58155),
    .O(net_58197)
  );
  ClkMux inmux_14_13_5_58207 (
    .I(net_5),
    .O(net_58207)
  );
  SRMux inmux_14_13_9_58208 (
    .I(net_9),
    .O(net_58208)
  );
  InMux inmux_14_14_58250_58319 (
    .I(net_58250),
    .O(net_58319)
  );
  InMux inmux_14_14_58251_58284 (
    .I(net_58251),
    .O(net_58284)
  );
  InMux inmux_14_14_58251_58296 (
    .I(net_58251),
    .O(net_58296)
  );
  InMux inmux_14_14_58251_58308 (
    .I(net_58251),
    .O(net_58308)
  );
  InMux inmux_14_14_58251_58313 (
    .I(net_58251),
    .O(net_58313)
  );
  InMux inmux_14_14_58251_58327 (
    .I(net_58251),
    .O(net_58327)
  );
  InMux inmux_14_14_58253_58322 (
    .I(net_58253),
    .O(net_58322)
  );
  InMux inmux_14_14_58254_58307 (
    .I(net_58254),
    .O(net_58307)
  );
  InMux inmux_14_14_58264_58320 (
    .I(net_58264),
    .O(net_58320)
  );
  InMux inmux_14_14_58268_58314 (
    .I(net_58268),
    .O(net_58314)
  );
  InMux inmux_14_14_58270_58285 (
    .I(net_58270),
    .O(net_58285)
  );
  InMux inmux_14_14_58273_58298 (
    .I(net_58273),
    .O(net_58298)
  );
  InMux inmux_14_14_58274_58325 (
    .I(net_58274),
    .O(net_58325)
  );
  InMux inmux_14_14_58275_58321 (
    .I(net_58275),
    .O(net_58321)
  );
  ClkMux inmux_14_14_5_58330 (
    .I(net_5),
    .O(net_58330)
  );
  CEMux inmux_14_14_6_58329 (
    .I(net_6),
    .O(net_58329)
  );
  SRMux inmux_14_14_9_58331 (
    .I(net_9),
    .O(net_58331)
  );
  InMux inmux_14_15_58373_58449 (
    .I(net_58373),
    .O(net_58449)
  );
  InMux inmux_14_15_58375_58427 (
    .I(net_58375),
    .O(net_58427)
  );
  InMux inmux_14_15_58378_58407 (
    .I(net_58378),
    .O(net_58407)
  );
  InMux inmux_14_15_58380_58419 (
    .I(net_58380),
    .O(net_58419)
  );
  InMux inmux_14_15_58385_58436 (
    .I(net_58385),
    .O(net_58436)
  );
  InMux inmux_14_15_58386_58415 (
    .I(net_58386),
    .O(net_58415)
  );
  InMux inmux_14_15_58387_58431 (
    .I(net_58387),
    .O(net_58431)
  );
  InMux inmux_14_15_58388_58444 (
    .I(net_58388),
    .O(net_58444)
  );
  InMux inmux_14_15_58393_58413 (
    .I(net_58393),
    .O(net_58413)
  );
  InMux inmux_14_15_58396_58412 (
    .I(net_58396),
    .O(net_58412)
  );
  ClkMux inmux_14_15_5_58453 (
    .I(net_5),
    .O(net_58453)
  );
  SRMux inmux_14_15_9_58454 (
    .I(net_9),
    .O(net_58454)
  );
  InMux inmux_14_16_58496_58567 (
    .I(net_58496),
    .O(net_58567)
  );
  InMux inmux_14_16_58499_58566 (
    .I(net_58499),
    .O(net_58566)
  );
  InMux inmux_14_16_58500_58572 (
    .I(net_58500),
    .O(net_58572)
  );
  InMux inmux_14_16_58501_58549 (
    .I(net_58501),
    .O(net_58549)
  );
  InMux inmux_14_16_58503_58542 (
    .I(net_58503),
    .O(net_58542)
  );
  InMux inmux_14_16_58504_58573 (
    .I(net_58504),
    .O(net_58573)
  );
  InMux inmux_14_16_58506_58554 (
    .I(net_58506),
    .O(net_58554)
  );
  InMux inmux_14_16_58507_58531 (
    .I(net_58507),
    .O(net_58531)
  );
  InMux inmux_14_16_58509_58543 (
    .I(net_58509),
    .O(net_58543)
  );
  InMux inmux_14_16_58510_58561 (
    .I(net_58510),
    .O(net_58561)
  );
  InMux inmux_14_16_58511_58555 (
    .I(net_58511),
    .O(net_58555)
  );
  InMux inmux_14_16_58514_58536 (
    .I(net_58514),
    .O(net_58536)
  );
  InMux inmux_14_16_58516_58560 (
    .I(net_58516),
    .O(net_58560)
  );
  InMux inmux_14_16_58522_58537 (
    .I(net_58522),
    .O(net_58537)
  );
  InMux inmux_14_16_58527_58548 (
    .I(net_58527),
    .O(net_58548)
  );
  InMux inmux_14_16_58534_58544 (
    .I(net_58534),
    .O(net_58544)
  );
  InMux inmux_14_16_58540_58550 (
    .I(net_58540),
    .O(net_58550)
  );
  InMux inmux_14_16_58546_58556 (
    .I(net_58546),
    .O(net_58556)
  );
  InMux inmux_14_16_58552_58562 (
    .I(net_58552),
    .O(net_58562)
  );
  InMux inmux_14_16_58558_58568 (
    .I(net_58558),
    .O(net_58568)
  );
  InMux inmux_14_16_58564_58574 (
    .I(net_58564),
    .O(net_58574)
  );
  ClkMux inmux_14_16_5_58576 (
    .I(net_5),
    .O(net_58576)
  );
  SRMux inmux_14_16_9_58577 (
    .I(net_9),
    .O(net_58577)
  );
  InMux inmux_14_17_58614_58655 (
    .I(net_58614),
    .O(net_58655)
  );
  InMux inmux_14_17_58620_58665 (
    .I(net_58620),
    .O(net_58665)
  );
  InMux inmux_14_17_58621_58685 (
    .I(net_58621),
    .O(net_58685)
  );
  InMux inmux_14_17_58621_58690 (
    .I(net_58621),
    .O(net_58690)
  );
  InMux inmux_14_17_58626_58653 (
    .I(net_58626),
    .O(net_58653)
  );
  InMux inmux_14_17_58630_58697 (
    .I(net_58630),
    .O(net_58697)
  );
  InMux inmux_14_17_58633_58672 (
    .I(net_58633),
    .O(net_58672)
  );
  InMux inmux_14_17_58646_58654 (
    .I(net_58646),
    .O(net_58654)
  );
  InMux inmux_14_17_58651_58661 (
    .I(net_58651),
    .O(net_58661)
  );
  ClkMux inmux_14_17_5_58699 (
    .I(net_5),
    .O(net_58699)
  );
  SRMux inmux_14_17_9_58700 (
    .I(net_9),
    .O(net_58700)
  );
  InMux inmux_14_18_58742_58775 (
    .I(net_58742),
    .O(net_58775)
  );
  InMux inmux_14_18_58743_58781 (
    .I(net_58743),
    .O(net_58781)
  );
  InMux inmux_14_18_58745_58795 (
    .I(net_58745),
    .O(net_58795)
  );
  InMux inmux_14_18_58747_58788 (
    .I(net_58747),
    .O(net_58788)
  );
  InMux inmux_14_18_58748_58794 (
    .I(net_58748),
    .O(net_58794)
  );
  InMux inmux_14_18_58750_58783 (
    .I(net_58750),
    .O(net_58783)
  );
  InMux inmux_14_18_58751_58789 (
    .I(net_58751),
    .O(net_58789)
  );
  InMux inmux_14_18_58751_58811 (
    .I(net_58751),
    .O(net_58811)
  );
  InMux inmux_14_18_58751_58818 (
    .I(net_58751),
    .O(net_58818)
  );
  InMux inmux_14_18_58752_58776 (
    .I(net_58752),
    .O(net_58776)
  );
  InMux inmux_14_18_58753_58777 (
    .I(net_58753),
    .O(net_58777)
  );
  InMux inmux_14_18_58753_58782 (
    .I(net_58753),
    .O(net_58782)
  );
  InMux inmux_14_18_58753_58787 (
    .I(net_58753),
    .O(net_58787)
  );
  InMux inmux_14_18_58753_58796 (
    .I(net_58753),
    .O(net_58796)
  );
  InMux inmux_14_18_58753_58808 (
    .I(net_58753),
    .O(net_58808)
  );
  InMux inmux_14_18_58753_58820 (
    .I(net_58753),
    .O(net_58820)
  );
  InMux inmux_14_18_58754_58817 (
    .I(net_58754),
    .O(net_58817)
  );
  InMux inmux_14_18_58756_58790 (
    .I(net_58756),
    .O(net_58790)
  );
  InMux inmux_14_18_58761_58807 (
    .I(net_58761),
    .O(net_58807)
  );
  InMux inmux_14_18_58764_58813 (
    .I(net_58764),
    .O(net_58813)
  );
  InMux inmux_14_18_58765_58814 (
    .I(net_58765),
    .O(net_58814)
  );
  InMux inmux_14_18_58768_58812 (
    .I(net_58768),
    .O(net_58812)
  );
  InMux inmux_14_18_58769_58806 (
    .I(net_58769),
    .O(net_58806)
  );
  InMux inmux_14_18_58770_58819 (
    .I(net_58770),
    .O(net_58819)
  );
  ClkMux inmux_14_18_5_58822 (
    .I(net_5),
    .O(net_58822)
  );
  CEMux inmux_14_18_6_58821 (
    .I(net_6),
    .O(net_58821)
  );
  SRMux inmux_14_18_9_58823 (
    .I(net_9),
    .O(net_58823)
  );
  CEMux inmux_14_19_58883_58944 (
    .I(net_58883),
    .O(net_58944)
  );
  InMux inmux_14_19_58884_58918 (
    .I(net_58884),
    .O(net_58918)
  );
  InMux inmux_14_19_58889_58916 (
    .I(net_58889),
    .O(net_58916)
  );
  InMux inmux_14_19_58892_58917 (
    .I(net_58892),
    .O(net_58917)
  );
  InMux inmux_14_19_58896_58919 (
    .I(net_58896),
    .O(net_58919)
  );
  ClkMux inmux_14_19_5_58945 (
    .I(net_5),
    .O(net_58945)
  );
  SRMux inmux_14_19_9_58946 (
    .I(net_9),
    .O(net_58946)
  );
  InMux inmux_14_1_56614_56683 (
    .I(net_56614),
    .O(net_56683)
  );
  InMux inmux_14_1_56627_56682 (
    .I(net_56627),
    .O(net_56682)
  );
  InMux inmux_14_2_56774_56826 (
    .I(net_56774),
    .O(net_56826)
  );
  InMux inmux_14_2_56776_56828 (
    .I(net_56776),
    .O(net_56828)
  );
  InMux inmux_14_2_56779_56820 (
    .I(net_56779),
    .O(net_56820)
  );
  InMux inmux_14_2_56783_56845 (
    .I(net_56783),
    .O(net_56845)
  );
  InMux inmux_14_2_56785_56809 (
    .I(net_56785),
    .O(net_56809)
  );
  InMux inmux_14_2_56788_56827 (
    .I(net_56788),
    .O(net_56827)
  );
  ClkMux inmux_14_2_5_56854 (
    .I(net_5),
    .O(net_56854)
  );
  CEMux inmux_14_2_8_56853 (
    .I(net_8),
    .O(net_56853)
  );
  SRMux inmux_14_2_9_56855 (
    .I(net_9),
    .O(net_56855)
  );
  InMux inmux_14_3_56900_56969 (
    .I(net_56900),
    .O(net_56969)
  );
  InMux inmux_14_3_56907_56972 (
    .I(net_56907),
    .O(net_56972)
  );
  ClkMux inmux_14_3_5_56977 (
    .I(net_5),
    .O(net_56977)
  );
  CEMux inmux_14_3_8_56976 (
    .I(net_8),
    .O(net_56976)
  );
  SRMux inmux_14_3_9_56978 (
    .I(net_9),
    .O(net_56978)
  );
  InMux inmux_14_4_57020_57096 (
    .I(net_57020),
    .O(net_57096)
  );
  InMux inmux_14_4_57026_57067 (
    .I(net_57026),
    .O(net_57067)
  );
  InMux inmux_14_4_57032_57071 (
    .I(net_57032),
    .O(net_57071)
  );
  InMux inmux_14_4_57035_57065 (
    .I(net_57035),
    .O(net_57065)
  );
  InMux inmux_14_4_57040_57079 (
    .I(net_57040),
    .O(net_57079)
  );
  InMux inmux_14_4_57043_57066 (
    .I(net_57043),
    .O(net_57066)
  );
  InMux inmux_14_4_57045_57089 (
    .I(net_57045),
    .O(net_57089)
  );
  InMux inmux_14_4_57048_57083 (
    .I(net_57048),
    .O(net_57083)
  );
  InMux inmux_14_4_57051_57055 (
    .I(net_57051),
    .O(net_57055)
  );
  ClkMux inmux_14_4_5_57100 (
    .I(net_5),
    .O(net_57100)
  );
  CEMux inmux_14_4_8_57099 (
    .I(net_8),
    .O(net_57099)
  );
  InMux inmux_14_5_57143_57207 (
    .I(net_57143),
    .O(net_57207)
  );
  InMux inmux_14_5_57145_57178 (
    .I(net_57145),
    .O(net_57178)
  );
  InMux inmux_14_5_57146_57179 (
    .I(net_57146),
    .O(net_57179)
  );
  InMux inmux_14_5_57152_57188 (
    .I(net_57152),
    .O(net_57188)
  );
  InMux inmux_14_5_57155_57218 (
    .I(net_57155),
    .O(net_57218)
  );
  InMux inmux_14_5_57156_57200 (
    .I(net_57156),
    .O(net_57200)
  );
  InMux inmux_14_5_57159_57183 (
    .I(net_57159),
    .O(net_57183)
  );
  InMux inmux_14_5_57160_57201 (
    .I(net_57160),
    .O(net_57201)
  );
  InMux inmux_14_5_57162_57177 (
    .I(net_57162),
    .O(net_57177)
  );
  InMux inmux_14_5_57162_57203 (
    .I(net_57162),
    .O(net_57203)
  );
  InMux inmux_14_5_57163_57197 (
    .I(net_57163),
    .O(net_57197)
  );
  InMux inmux_14_5_57165_57202 (
    .I(net_57165),
    .O(net_57202)
  );
  InMux inmux_14_5_57166_57208 (
    .I(net_57166),
    .O(net_57208)
  );
  InMux inmux_14_5_57168_57214 (
    .I(net_57168),
    .O(net_57214)
  );
  CEMux inmux_14_5_57170_57222 (
    .I(net_57170),
    .O(net_57222)
  );
  InMux inmux_14_5_57172_57209 (
    .I(net_57172),
    .O(net_57209)
  );
  InMux inmux_14_5_57173_57206 (
    .I(net_57173),
    .O(net_57206)
  );
  InMux inmux_14_5_57174_57176 (
    .I(net_57174),
    .O(net_57176)
  );
  ClkMux inmux_14_5_5_57223 (
    .I(net_5),
    .O(net_57223)
  );
  InMux inmux_14_6_57266_57337 (
    .I(net_57266),
    .O(net_57337)
  );
  InMux inmux_14_6_57269_57319 (
    .I(net_57269),
    .O(net_57319)
  );
  InMux inmux_14_6_57270_57325 (
    .I(net_57270),
    .O(net_57325)
  );
  InMux inmux_14_6_57273_57341 (
    .I(net_57273),
    .O(net_57341)
  );
  InMux inmux_14_6_57275_57344 (
    .I(net_57275),
    .O(net_57344)
  );
  InMux inmux_14_6_57276_57317 (
    .I(net_57276),
    .O(net_57317)
  );
  InMux inmux_14_6_57277_57308 (
    .I(net_57277),
    .O(net_57308)
  );
  InMux inmux_14_6_57277_57342 (
    .I(net_57277),
    .O(net_57342)
  );
  InMux inmux_14_6_57278_57326 (
    .I(net_57278),
    .O(net_57326)
  );
  InMux inmux_14_6_57279_57320 (
    .I(net_57279),
    .O(net_57320)
  );
  InMux inmux_14_6_57282_57332 (
    .I(net_57282),
    .O(net_57332)
  );
  InMux inmux_14_6_57288_57318 (
    .I(net_57288),
    .O(net_57318)
  );
  InMux inmux_14_6_57290_57307 (
    .I(net_57290),
    .O(net_57307)
  );
  InMux inmux_14_6_57294_57302 (
    .I(net_57294),
    .O(net_57302)
  );
  InMux inmux_14_6_57295_57306 (
    .I(net_57295),
    .O(net_57306)
  );
  InMux inmux_14_6_57296_57305 (
    .I(net_57296),
    .O(net_57305)
  );
  InMux inmux_14_6_57296_57343 (
    .I(net_57296),
    .O(net_57343)
  );
  ClkMux inmux_14_6_5_57346 (
    .I(net_5),
    .O(net_57346)
  );
  SRMux inmux_14_6_9_57347 (
    .I(net_9),
    .O(net_57347)
  );
  InMux inmux_14_7_57396_57440 (
    .I(net_57396),
    .O(net_57440)
  );
  InMux inmux_14_7_57402_57465 (
    .I(net_57402),
    .O(net_57465)
  );
  InMux inmux_14_7_57404_57460 (
    .I(net_57404),
    .O(net_57460)
  );
  InMux inmux_14_7_57407_57429 (
    .I(net_57407),
    .O(net_57429)
  );
  InMux inmux_14_7_57416_57455 (
    .I(net_57416),
    .O(net_57455)
  );
  ClkMux inmux_14_7_5_57469 (
    .I(net_5),
    .O(net_57469)
  );
  SRMux inmux_14_7_9_57470 (
    .I(net_9),
    .O(net_57470)
  );
  InMux inmux_14_8_57512_57583 (
    .I(net_57512),
    .O(net_57583)
  );
  InMux inmux_14_8_57513_57587 (
    .I(net_57513),
    .O(net_57587)
  );
  InMux inmux_14_8_57517_57584 (
    .I(net_57517),
    .O(net_57584)
  );
  InMux inmux_14_8_57521_57547 (
    .I(net_57521),
    .O(net_57547)
  );
  InMux inmux_14_8_57523_57559 (
    .I(net_57523),
    .O(net_57559)
  );
  InMux inmux_14_8_57524_57570 (
    .I(net_57524),
    .O(net_57570)
  );
  InMux inmux_14_8_57525_57552 (
    .I(net_57525),
    .O(net_57552)
  );
  InMux inmux_14_8_57528_57576 (
    .I(net_57528),
    .O(net_57576)
  );
  InMux inmux_14_8_57536_57582 (
    .I(net_57536),
    .O(net_57582)
  );
  InMux inmux_14_8_57538_57563 (
    .I(net_57538),
    .O(net_57563)
  );
  InMux inmux_14_8_57541_57581 (
    .I(net_57541),
    .O(net_57581)
  );
  ClkMux inmux_14_8_5_57592 (
    .I(net_5),
    .O(net_57592)
  );
  SRMux inmux_14_8_9_57593 (
    .I(net_9),
    .O(net_57593)
  );
  InMux inmux_14_9_57635_57706 (
    .I(net_57635),
    .O(net_57706)
  );
  InMux inmux_14_9_57636_57705 (
    .I(net_57636),
    .O(net_57705)
  );
  InMux inmux_14_9_57637_57675 (
    .I(net_57637),
    .O(net_57675)
  );
  InMux inmux_14_9_57639_57668 (
    .I(net_57639),
    .O(net_57668)
  );
  InMux inmux_14_9_57643_57707 (
    .I(net_57643),
    .O(net_57707)
  );
  InMux inmux_14_9_57644_57704 (
    .I(net_57644),
    .O(net_57704)
  );
  CEMux inmux_14_9_57646_57714 (
    .I(net_57646),
    .O(net_57714)
  );
  ClkMux inmux_14_9_5_57715 (
    .I(net_5),
    .O(net_57715)
  );
  ClkMux inmux_15_10_5_61668 (
    .I(net_5),
    .O(net_61668)
  );
  InMux inmux_15_10_61588_61633 (
    .I(net_61588),
    .O(net_61633)
  );
  InMux inmux_15_10_61588_61664 (
    .I(net_61588),
    .O(net_61664)
  );
  InMux inmux_15_10_61594_61666 (
    .I(net_61594),
    .O(net_61666)
  );
  InMux inmux_15_10_61596_61627 (
    .I(net_61596),
    .O(net_61627)
  );
  InMux inmux_15_10_61596_61641 (
    .I(net_61596),
    .O(net_61641)
  );
  InMux inmux_15_10_61597_61628 (
    .I(net_61597),
    .O(net_61628)
  );
  InMux inmux_15_10_61602_61622 (
    .I(net_61602),
    .O(net_61622)
  );
  CEMux inmux_15_10_61606_61667 (
    .I(net_61606),
    .O(net_61667)
  );
  InMux inmux_15_10_61607_61639 (
    .I(net_61607),
    .O(net_61639)
  );
  InMux inmux_15_10_61610_61630 (
    .I(net_61610),
    .O(net_61630)
  );
  InMux inmux_15_10_61610_61657 (
    .I(net_61610),
    .O(net_61657)
  );
  InMux inmux_15_10_61614_61634 (
    .I(net_61614),
    .O(net_61634)
  );
  InMux inmux_15_10_61626_61636 (
    .I(net_61626),
    .O(net_61636)
  );
  InMux inmux_15_10_61632_61642 (
    .I(net_61632),
    .O(net_61642)
  );
  SRMux inmux_15_10_9_61669 (
    .I(net_9),
    .O(net_61669)
  );
  ClkMux inmux_15_11_5_61791 (
    .I(net_5),
    .O(net_61791)
  );
  InMux inmux_15_11_61713_61753 (
    .I(net_61713),
    .O(net_61753)
  );
  InMux inmux_15_11_61714_61752 (
    .I(net_61714),
    .O(net_61752)
  );
  InMux inmux_15_11_61720_61746 (
    .I(net_61720),
    .O(net_61746)
  );
  InMux inmux_15_11_61723_61776 (
    .I(net_61723),
    .O(net_61776)
  );
  InMux inmux_15_11_61724_61780 (
    .I(net_61724),
    .O(net_61780)
  );
  InMux inmux_15_11_61725_61747 (
    .I(net_61725),
    .O(net_61747)
  );
  InMux inmux_15_11_61731_61765 (
    .I(net_61731),
    .O(net_61765)
  );
  InMux inmux_15_11_61733_61756 (
    .I(net_61733),
    .O(net_61756)
  );
  InMux inmux_15_11_61734_61788 (
    .I(net_61734),
    .O(net_61788)
  );
  InMux inmux_15_11_61736_61744 (
    .I(net_61736),
    .O(net_61744)
  );
  InMux inmux_15_11_61737_61769 (
    .I(net_61737),
    .O(net_61769)
  );
  InMux inmux_15_11_61742_61751 (
    .I(net_61742),
    .O(net_61751)
  );
  SRMux inmux_15_11_9_61792 (
    .I(net_9),
    .O(net_61792)
  );
  ClkMux inmux_15_12_5_61914 (
    .I(net_5),
    .O(net_61914)
  );
  InMux inmux_15_12_61841_61887 (
    .I(net_61841),
    .O(net_61887)
  );
  InMux inmux_15_12_61843_61891 (
    .I(net_61843),
    .O(net_61891)
  );
  InMux inmux_15_12_61849_61903 (
    .I(net_61849),
    .O(net_61903)
  );
  InMux inmux_15_12_61851_61899 (
    .I(net_61851),
    .O(net_61899)
  );
  InMux inmux_15_12_61852_61869 (
    .I(net_61852),
    .O(net_61869)
  );
  InMux inmux_15_12_61854_61874 (
    .I(net_61854),
    .O(net_61874)
  );
  InMux inmux_15_12_61857_61882 (
    .I(net_61857),
    .O(net_61882)
  );
  InMux inmux_15_12_61864_61870 (
    .I(net_61864),
    .O(net_61870)
  );
  InMux inmux_15_12_61865_61910 (
    .I(net_61865),
    .O(net_61910)
  );
  SRMux inmux_15_12_9_61915 (
    .I(net_9),
    .O(net_61915)
  );
  ClkMux inmux_15_13_5_62037 (
    .I(net_5),
    .O(net_62037)
  );
  InMux inmux_15_13_61962_61991 (
    .I(net_61962),
    .O(net_61991)
  );
  InMux inmux_15_13_61968_61992 (
    .I(net_61968),
    .O(net_61992)
  );
  InMux inmux_15_13_61975_62004 (
    .I(net_61975),
    .O(net_62004)
  );
  InMux inmux_15_13_61976_62010 (
    .I(net_61976),
    .O(net_62010)
  );
  InMux inmux_15_13_61982_61997 (
    .I(net_61982),
    .O(net_61997)
  );
  InMux inmux_15_13_61985_62015 (
    .I(net_61985),
    .O(net_62015)
  );
  InMux inmux_15_13_61986_62021 (
    .I(net_61986),
    .O(net_62021)
  );
  InMux inmux_15_13_61987_62027 (
    .I(net_61987),
    .O(net_62027)
  );
  InMux inmux_15_13_61989_61999 (
    .I(net_61989),
    .O(net_61999)
  );
  InMux inmux_15_13_61995_62005 (
    .I(net_61995),
    .O(net_62005)
  );
  InMux inmux_15_13_62001_62011 (
    .I(net_62001),
    .O(net_62011)
  );
  InMux inmux_15_13_62007_62017 (
    .I(net_62007),
    .O(net_62017)
  );
  InMux inmux_15_13_62013_62023 (
    .I(net_62013),
    .O(net_62023)
  );
  InMux inmux_15_13_62019_62029 (
    .I(net_62019),
    .O(net_62029)
  );
  InMux inmux_15_13_62025_62035 (
    .I(net_62025),
    .O(net_62035)
  );
  SRMux inmux_15_13_9_62038 (
    .I(net_9),
    .O(net_62038)
  );
  ClkMux inmux_15_14_5_62160 (
    .I(net_5),
    .O(net_62160)
  );
  InMux inmux_15_14_62081_62138 (
    .I(net_62081),
    .O(net_62138)
  );
  InMux inmux_15_14_62082_62127 (
    .I(net_62082),
    .O(net_62127)
  );
  InMux inmux_15_14_62083_62150 (
    .I(net_62083),
    .O(net_62150)
  );
  InMux inmux_15_14_62085_62131 (
    .I(net_62085),
    .O(net_62131)
  );
  InMux inmux_15_14_62090_62121 (
    .I(net_62090),
    .O(net_62121)
  );
  InMux inmux_15_14_62090_62128 (
    .I(net_62090),
    .O(net_62128)
  );
  InMux inmux_15_14_62090_62133 (
    .I(net_62090),
    .O(net_62133)
  );
  InMux inmux_15_14_62090_62140 (
    .I(net_62090),
    .O(net_62140)
  );
  InMux inmux_15_14_62090_62152 (
    .I(net_62090),
    .O(net_62152)
  );
  CEMux inmux_15_14_62091_62159 (
    .I(net_62091),
    .O(net_62159)
  );
  InMux inmux_15_14_62092_62145 (
    .I(net_62092),
    .O(net_62145)
  );
  InMux inmux_15_14_62093_62156 (
    .I(net_62093),
    .O(net_62156)
  );
  InMux inmux_15_14_62096_62144 (
    .I(net_62096),
    .O(net_62144)
  );
  InMux inmux_15_14_62097_62119 (
    .I(net_62097),
    .O(net_62119)
  );
  InMux inmux_15_14_62107_62158 (
    .I(net_62107),
    .O(net_62158)
  );
  InMux inmux_15_14_62109_62115 (
    .I(net_62109),
    .O(net_62115)
  );
  SRMux inmux_15_14_9_62161 (
    .I(net_9),
    .O(net_62161)
  );
  ClkMux inmux_15_15_5_62283 (
    .I(net_5),
    .O(net_62283)
  );
  InMux inmux_15_15_62212_62250 (
    .I(net_62212),
    .O(net_62250)
  );
  InMux inmux_15_15_62213_62261 (
    .I(net_62213),
    .O(net_62261)
  );
  InMux inmux_15_15_62214_62236 (
    .I(net_62214),
    .O(net_62236)
  );
  InMux inmux_15_15_62228_62272 (
    .I(net_62228),
    .O(net_62272)
  );
  InMux inmux_15_15_62232_62245 (
    .I(net_62232),
    .O(net_62245)
  );
  InMux inmux_15_15_62233_62256 (
    .I(net_62233),
    .O(net_62256)
  );
  InMux inmux_15_15_62233_62280 (
    .I(net_62233),
    .O(net_62280)
  );
  SRMux inmux_15_15_9_62284 (
    .I(net_9),
    .O(net_62284)
  );
  ClkMux inmux_15_16_5_62406 (
    .I(net_5),
    .O(net_62406)
  );
  InMux inmux_15_16_62326_62366 (
    .I(net_62326),
    .O(net_62366)
  );
  InMux inmux_15_16_62327_62384 (
    .I(net_62327),
    .O(net_62384)
  );
  InMux inmux_15_16_62331_62396 (
    .I(net_62331),
    .O(net_62396)
  );
  InMux inmux_15_16_62333_62391 (
    .I(net_62333),
    .O(net_62391)
  );
  InMux inmux_15_16_62335_62378 (
    .I(net_62335),
    .O(net_62378)
  );
  InMux inmux_15_16_62337_62402 (
    .I(net_62337),
    .O(net_62402)
  );
  InMux inmux_15_16_62342_62397 (
    .I(net_62342),
    .O(net_62397)
  );
  InMux inmux_15_16_62345_62367 (
    .I(net_62345),
    .O(net_62367)
  );
  InMux inmux_15_16_62347_62372 (
    .I(net_62347),
    .O(net_62372)
  );
  InMux inmux_15_16_62348_62373 (
    .I(net_62348),
    .O(net_62373)
  );
  InMux inmux_15_16_62351_62385 (
    .I(net_62351),
    .O(net_62385)
  );
  InMux inmux_15_16_62352_62379 (
    .I(net_62352),
    .O(net_62379)
  );
  InMux inmux_15_16_62353_62361 (
    .I(net_62353),
    .O(net_62361)
  );
  InMux inmux_15_16_62353_62368 (
    .I(net_62353),
    .O(net_62368)
  );
  InMux inmux_15_16_62355_62390 (
    .I(net_62355),
    .O(net_62390)
  );
  InMux inmux_15_16_62356_62403 (
    .I(net_62356),
    .O(net_62403)
  );
  InMux inmux_15_16_62364_62374 (
    .I(net_62364),
    .O(net_62374)
  );
  InMux inmux_15_16_62370_62380 (
    .I(net_62370),
    .O(net_62380)
  );
  InMux inmux_15_16_62376_62386 (
    .I(net_62376),
    .O(net_62386)
  );
  InMux inmux_15_16_62382_62392 (
    .I(net_62382),
    .O(net_62392)
  );
  InMux inmux_15_16_62388_62398 (
    .I(net_62388),
    .O(net_62398)
  );
  InMux inmux_15_16_62394_62404 (
    .I(net_62394),
    .O(net_62404)
  );
  SRMux inmux_15_16_9_62407 (
    .I(net_9),
    .O(net_62407)
  );
  ClkMux inmux_15_17_5_62529 (
    .I(net_5),
    .O(net_62529)
  );
  InMux inmux_15_17_62444_62485 (
    .I(net_62444),
    .O(net_62485)
  );
  InMux inmux_15_17_62449_62496 (
    .I(net_62449),
    .O(net_62496)
  );
  InMux inmux_15_17_62466_62509 (
    .I(net_62466),
    .O(net_62509)
  );
  InMux inmux_15_17_62467_62506 (
    .I(net_62467),
    .O(net_62506)
  );
  InMux inmux_15_17_62468_62483 (
    .I(net_62468),
    .O(net_62483)
  );
  InMux inmux_15_17_62470_62507 (
    .I(net_62470),
    .O(net_62507)
  );
  InMux inmux_15_17_62480_62484 (
    .I(net_62480),
    .O(net_62484)
  );
  InMux inmux_15_17_62481_62491 (
    .I(net_62481),
    .O(net_62491)
  );
  SRMux inmux_15_17_9_62530 (
    .I(net_9),
    .O(net_62530)
  );
  ClkMux inmux_15_18_5_62652 (
    .I(net_5),
    .O(net_62652)
  );
  InMux inmux_15_18_62575_62632 (
    .I(net_62575),
    .O(net_62632)
  );
  InMux inmux_15_18_62582_62630 (
    .I(net_62582),
    .O(net_62630)
  );
  CEMux inmux_15_18_62583_62651 (
    .I(net_62583),
    .O(net_62651)
  );
  InMux inmux_15_18_62592_62629 (
    .I(net_62592),
    .O(net_62629)
  );
  InMux inmux_15_18_62597_62631 (
    .I(net_62597),
    .O(net_62631)
  );
  SRMux inmux_15_18_9_62653 (
    .I(net_9),
    .O(net_62653)
  );
  CEMux inmux_15_2_12_60683 (
    .I(net_12),
    .O(net_60683)
  );
  ClkMux inmux_15_2_5_60684 (
    .I(net_5),
    .O(net_60684)
  );
  InMux inmux_15_2_60627_60676 (
    .I(net_60627),
    .O(net_60676)
  );
  ClkMux inmux_15_3_5_60807 (
    .I(net_5),
    .O(net_60807)
  );
  InMux inmux_15_3_60729_60784 (
    .I(net_60729),
    .O(net_60784)
  );
  InMux inmux_15_3_60731_60774 (
    .I(net_60731),
    .O(net_60774)
  );
  SRMux inmux_15_3_9_60808 (
    .I(net_9),
    .O(net_60808)
  );
  ClkMux inmux_15_4_5_60930 (
    .I(net_5),
    .O(net_60930)
  );
  InMux inmux_15_4_60850_60926 (
    .I(net_60850),
    .O(net_60926)
  );
  InMux inmux_15_4_60852_60890 (
    .I(net_60852),
    .O(net_60890)
  );
  InMux inmux_15_4_60852_60904 (
    .I(net_60852),
    .O(net_60904)
  );
  InMux inmux_15_4_60852_60909 (
    .I(net_60852),
    .O(net_60909)
  );
  InMux inmux_15_4_60852_60914 (
    .I(net_60852),
    .O(net_60914)
  );
  InMux inmux_15_4_60852_60921 (
    .I(net_60852),
    .O(net_60921)
  );
  InMux inmux_15_4_60860_60901 (
    .I(net_60860),
    .O(net_60901)
  );
  InMux inmux_15_4_60866_60892 (
    .I(net_60866),
    .O(net_60892)
  );
  InMux inmux_15_4_60870_60895 (
    .I(net_60870),
    .O(net_60895)
  );
  InMux inmux_15_4_60874_60908 (
    .I(net_60874),
    .O(net_60908)
  );
  InMux inmux_15_4_60876_60922 (
    .I(net_60876),
    .O(net_60922)
  );
  InMux inmux_15_4_60878_60915 (
    .I(net_60878),
    .O(net_60915)
  );
  InMux inmux_15_4_60880_60886 (
    .I(net_60880),
    .O(net_60886)
  );
  SRMux inmux_15_4_9_60931 (
    .I(net_9),
    .O(net_60931)
  );
  ClkMux inmux_15_5_5_61053 (
    .I(net_5),
    .O(net_61053)
  );
  InMux inmux_15_5_60973_61020 (
    .I(net_60973),
    .O(net_61020)
  );
  InMux inmux_15_5_60978_61033 (
    .I(net_60978),
    .O(net_61033)
  );
  InMux inmux_15_5_60982_61025 (
    .I(net_60982),
    .O(net_61025)
  );
  InMux inmux_15_5_60983_61036 (
    .I(net_60983),
    .O(net_61036)
  );
  InMux inmux_15_5_60988_61042 (
    .I(net_60988),
    .O(net_61042)
  );
  InMux inmux_15_5_60991_61006 (
    .I(net_60991),
    .O(net_61006)
  );
  InMux inmux_15_5_60991_61015 (
    .I(net_60991),
    .O(net_61015)
  );
  InMux inmux_15_5_60991_61018 (
    .I(net_60991),
    .O(net_61018)
  );
  InMux inmux_15_5_60991_61027 (
    .I(net_60991),
    .O(net_61027)
  );
  InMux inmux_15_5_60991_61032 (
    .I(net_60991),
    .O(net_61032)
  );
  InMux inmux_15_5_60991_61039 (
    .I(net_60991),
    .O(net_61039)
  );
  InMux inmux_15_5_60991_61044 (
    .I(net_60991),
    .O(net_61044)
  );
  InMux inmux_15_5_60991_61049 (
    .I(net_60991),
    .O(net_61049)
  );
  InMux inmux_15_5_60993_61051 (
    .I(net_60993),
    .O(net_61051)
  );
  InMux inmux_15_5_60998_61013 (
    .I(net_60998),
    .O(net_61013)
  );
  InMux inmux_15_5_61001_61007 (
    .I(net_61001),
    .O(net_61007)
  );
  SRMux inmux_15_5_9_61054 (
    .I(net_9),
    .O(net_61054)
  );
  ClkMux inmux_15_6_5_61176 (
    .I(net_5),
    .O(net_61176)
  );
  InMux inmux_15_6_61096_61129 (
    .I(net_61096),
    .O(net_61129)
  );
  InMux inmux_15_6_61097_61173 (
    .I(net_61097),
    .O(net_61173)
  );
  InMux inmux_15_6_61098_61148 (
    .I(net_61098),
    .O(net_61148)
  );
  InMux inmux_15_6_61099_61159 (
    .I(net_61099),
    .O(net_61159)
  );
  InMux inmux_15_6_61100_61174 (
    .I(net_61100),
    .O(net_61174)
  );
  InMux inmux_15_6_61102_61155 (
    .I(net_61102),
    .O(net_61155)
  );
  InMux inmux_15_6_61104_61147 (
    .I(net_61104),
    .O(net_61147)
  );
  InMux inmux_15_6_61106_61168 (
    .I(net_61106),
    .O(net_61168)
  );
  InMux inmux_15_6_61107_61165 (
    .I(net_61107),
    .O(net_61165)
  );
  InMux inmux_15_6_61108_61130 (
    .I(net_61108),
    .O(net_61130)
  );
  InMux inmux_15_6_61109_61162 (
    .I(net_61109),
    .O(net_61162)
  );
  InMux inmux_15_6_61111_61131 (
    .I(net_61111),
    .O(net_61131)
  );
  InMux inmux_15_6_61112_61172 (
    .I(net_61112),
    .O(net_61172)
  );
  InMux inmux_15_6_61114_61136 (
    .I(net_61114),
    .O(net_61136)
  );
  InMux inmux_15_6_61115_61154 (
    .I(net_61115),
    .O(net_61154)
  );
  InMux inmux_15_6_61116_61153 (
    .I(net_61116),
    .O(net_61153)
  );
  InMux inmux_15_6_61117_61135 (
    .I(net_61117),
    .O(net_61135)
  );
  InMux inmux_15_6_61118_61160 (
    .I(net_61118),
    .O(net_61160)
  );
  InMux inmux_15_6_61121_61150 (
    .I(net_61121),
    .O(net_61150)
  );
  InMux inmux_15_6_61122_61132 (
    .I(net_61122),
    .O(net_61132)
  );
  InMux inmux_15_6_61122_61137 (
    .I(net_61122),
    .O(net_61137)
  );
  InMux inmux_15_6_61122_61149 (
    .I(net_61122),
    .O(net_61149)
  );
  InMux inmux_15_6_61122_61161 (
    .I(net_61122),
    .O(net_61161)
  );
  InMux inmux_15_6_61122_61166 (
    .I(net_61122),
    .O(net_61166)
  );
  InMux inmux_15_6_61122_61171 (
    .I(net_61122),
    .O(net_61171)
  );
  CEMux inmux_15_6_61123_61175 (
    .I(net_61123),
    .O(net_61175)
  );
  InMux inmux_15_6_61124_61156 (
    .I(net_61124),
    .O(net_61156)
  );
  InMux inmux_15_6_61125_61138 (
    .I(net_61125),
    .O(net_61138)
  );
  InMux inmux_15_6_61127_61167 (
    .I(net_61127),
    .O(net_61167)
  );
  SRMux inmux_15_6_9_61177 (
    .I(net_9),
    .O(net_61177)
  );
  ClkMux inmux_15_7_5_61299 (
    .I(net_5),
    .O(net_61299)
  );
  InMux inmux_15_7_61234_61266 (
    .I(net_61234),
    .O(net_61266)
  );
  InMux inmux_15_7_61241_61276 (
    .I(net_61241),
    .O(net_61276)
  );
  InMux inmux_15_7_61242_61272 (
    .I(net_61242),
    .O(net_61272)
  );
  InMux inmux_15_7_61246_61290 (
    .I(net_61246),
    .O(net_61290)
  );
  SRMux inmux_15_7_9_61300 (
    .I(net_9),
    .O(net_61300)
  );
  ClkMux inmux_15_8_5_61422 (
    .I(net_5),
    .O(net_61422)
  );
  InMux inmux_15_8_61345_61390 (
    .I(net_61345),
    .O(net_61390)
  );
  InMux inmux_15_8_61347_61395 (
    .I(net_61347),
    .O(net_61395)
  );
  InMux inmux_15_8_61355_61382 (
    .I(net_61355),
    .O(net_61382)
  );
  InMux inmux_15_8_61366_61400 (
    .I(net_61366),
    .O(net_61400)
  );
  SRMux inmux_15_8_9_61423 (
    .I(net_9),
    .O(net_61423)
  );
  ClkMux inmux_15_9_5_61545 (
    .I(net_5),
    .O(net_61545)
  );
  InMux inmux_15_9_61468_61506 (
    .I(net_61468),
    .O(net_61506)
  );
  InMux inmux_15_9_61469_61498 (
    .I(net_61469),
    .O(net_61498)
  );
  InMux inmux_15_9_61475_61513 (
    .I(net_61475),
    .O(net_61513)
  );
  InMux inmux_15_9_61476_61536 (
    .I(net_61476),
    .O(net_61536)
  );
  InMux inmux_15_9_61485_61524 (
    .I(net_61485),
    .O(net_61524)
  );
  CEMux inmux_15_9_61492_61544 (
    .I(net_61492),
    .O(net_61544)
  );
  InMux inmux_15_9_61496_61519 (
    .I(net_61496),
    .O(net_61519)
  );
  IoInMux inmux_16_0_64225_64205 (
    .I(net_64225),
    .O(net_64205)
  );
  ClkMux inmux_16_10_5_65499 (
    .I(net_5),
    .O(net_65499)
  );
  InMux inmux_16_10_65421_65464 (
    .I(net_65421),
    .O(net_65464)
  );
  InMux inmux_16_10_65423_65478 (
    .I(net_65423),
    .O(net_65478)
  );
  InMux inmux_16_10_65427_65455 (
    .I(net_65427),
    .O(net_65455)
  );
  InMux inmux_16_10_65427_65465 (
    .I(net_65427),
    .O(net_65465)
  );
  InMux inmux_16_10_65427_65472 (
    .I(net_65427),
    .O(net_65472)
  );
  InMux inmux_16_10_65427_65477 (
    .I(net_65427),
    .O(net_65477)
  );
  InMux inmux_16_10_65427_65482 (
    .I(net_65427),
    .O(net_65482)
  );
  InMux inmux_16_10_65427_65489 (
    .I(net_65427),
    .O(net_65489)
  );
  InMux inmux_16_10_65427_65494 (
    .I(net_65427),
    .O(net_65494)
  );
  InMux inmux_16_10_65428_65454 (
    .I(net_65428),
    .O(net_65454)
  );
  InMux inmux_16_10_65436_65458 (
    .I(net_65436),
    .O(net_65458)
  );
  InMux inmux_16_10_65438_65491 (
    .I(net_65438),
    .O(net_65491)
  );
  InMux inmux_16_10_65439_65485 (
    .I(net_65439),
    .O(net_65485)
  );
  InMux inmux_16_10_65444_65495 (
    .I(net_65444),
    .O(net_65495)
  );
  InMux inmux_16_10_65445_65470 (
    .I(net_65445),
    .O(net_65470)
  );
  InMux inmux_16_10_65446_65461 (
    .I(net_65446),
    .O(net_65461)
  );
  SRMux inmux_16_10_9_65500 (
    .I(net_9),
    .O(net_65500)
  );
  ClkMux inmux_16_11_5_65622 (
    .I(net_5),
    .O(net_65622)
  );
  InMux inmux_16_11_65543_65576 (
    .I(net_65543),
    .O(net_65576)
  );
  InMux inmux_16_11_65543_65612 (
    .I(net_65543),
    .O(net_65612)
  );
  CEMux inmux_16_11_65544_65621 (
    .I(net_65544),
    .O(net_65621)
  );
  InMux inmux_16_11_65546_65577 (
    .I(net_65546),
    .O(net_65577)
  );
  InMux inmux_16_11_65546_65611 (
    .I(net_65546),
    .O(net_65611)
  );
  InMux inmux_16_11_65547_65595 (
    .I(net_65547),
    .O(net_65595)
  );
  InMux inmux_16_11_65547_65600 (
    .I(net_65547),
    .O(net_65600)
  );
  InMux inmux_16_11_65555_65589 (
    .I(net_65555),
    .O(net_65589)
  );
  InMux inmux_16_11_65562_65601 (
    .I(net_65562),
    .O(net_65601)
  );
  InMux inmux_16_11_65565_65581 (
    .I(net_65565),
    .O(net_65581)
  );
  InMux inmux_16_11_65565_65593 (
    .I(net_65565),
    .O(net_65593)
  );
  InMux inmux_16_11_65567_65582 (
    .I(net_65567),
    .O(net_65582)
  );
  InMux inmux_16_11_65568_65588 (
    .I(net_65568),
    .O(net_65588)
  );
  InMux inmux_16_11_65569_65594 (
    .I(net_65569),
    .O(net_65594)
  );
  InMux inmux_16_11_65571_65620 (
    .I(net_65571),
    .O(net_65620)
  );
  InMux inmux_16_11_65572_65583 (
    .I(net_65572),
    .O(net_65583)
  );
  InMux inmux_16_11_65573_65587 (
    .I(net_65573),
    .O(net_65587)
  );
  InMux inmux_16_11_65573_65599 (
    .I(net_65573),
    .O(net_65599)
  );
  InMux inmux_16_11_65573_65613 (
    .I(net_65573),
    .O(net_65613)
  );
  InMux inmux_16_11_65573_65618 (
    .I(net_65573),
    .O(net_65618)
  );
  InMux inmux_16_11_65574_65584 (
    .I(net_65574),
    .O(net_65584)
  );
  InMux inmux_16_11_65580_65590 (
    .I(net_65580),
    .O(net_65590)
  );
  InMux inmux_16_11_65586_65596 (
    .I(net_65586),
    .O(net_65596)
  );
  InMux inmux_16_11_65592_65602 (
    .I(net_65592),
    .O(net_65602)
  );
  InMux inmux_16_11_65598_65608 (
    .I(net_65598),
    .O(net_65608)
  );
  SRMux inmux_16_11_9_65623 (
    .I(net_9),
    .O(net_65623)
  );
  ClkMux inmux_16_12_5_65745 (
    .I(net_5),
    .O(net_65745)
  );
  CEMux inmux_16_12_65667_65744 (
    .I(net_65667),
    .O(net_65744)
  );
  InMux inmux_16_12_65668_65711 (
    .I(net_65668),
    .O(net_65711)
  );
  InMux inmux_16_12_65670_65713 (
    .I(net_65670),
    .O(net_65713)
  );
  InMux inmux_16_12_65672_65716 (
    .I(net_65672),
    .O(net_65716)
  );
  InMux inmux_16_12_65673_65718 (
    .I(net_65673),
    .O(net_65718)
  );
  InMux inmux_16_12_65674_65719 (
    .I(net_65674),
    .O(net_65719)
  );
  InMux inmux_16_12_65677_65735 (
    .I(net_65677),
    .O(net_65735)
  );
  InMux inmux_16_12_65678_65712 (
    .I(net_65678),
    .O(net_65712)
  );
  InMux inmux_16_12_65678_65717 (
    .I(net_65678),
    .O(net_65717)
  );
  InMux inmux_16_12_65678_65734 (
    .I(net_65678),
    .O(net_65734)
  );
  InMux inmux_16_12_65678_65741 (
    .I(net_65678),
    .O(net_65741)
  );
  InMux inmux_16_12_65679_65742 (
    .I(net_65679),
    .O(net_65742)
  );
  InMux inmux_16_12_65680_65743 (
    .I(net_65680),
    .O(net_65743)
  );
  InMux inmux_16_12_65682_65740 (
    .I(net_65682),
    .O(net_65740)
  );
  InMux inmux_16_12_65686_65737 (
    .I(net_65686),
    .O(net_65737)
  );
  InMux inmux_16_12_65690_65710 (
    .I(net_65690),
    .O(net_65710)
  );
  InMux inmux_16_12_65694_65736 (
    .I(net_65694),
    .O(net_65736)
  );
  ClkMux inmux_16_13_5_65868 (
    .I(net_5),
    .O(net_65868)
  );
  InMux inmux_16_13_65790_65847 (
    .I(net_65790),
    .O(net_65847)
  );
  InMux inmux_16_13_65792_65835 (
    .I(net_65792),
    .O(net_65835)
  );
  InMux inmux_16_13_65796_65834 (
    .I(net_65796),
    .O(net_65834)
  );
  InMux inmux_16_13_65797_65864 (
    .I(net_65797),
    .O(net_65864)
  );
  CEMux inmux_16_13_65799_65867 (
    .I(net_65799),
    .O(net_65867)
  );
  InMux inmux_16_13_65800_65829 (
    .I(net_65800),
    .O(net_65829)
  );
  InMux inmux_16_13_65806_65828 (
    .I(net_65806),
    .O(net_65828)
  );
  InMux inmux_16_13_65807_65846 (
    .I(net_65807),
    .O(net_65846)
  );
  InMux inmux_16_13_65810_65840 (
    .I(net_65810),
    .O(net_65840)
  );
  InMux inmux_16_13_65812_65822 (
    .I(net_65812),
    .O(net_65822)
  );
  InMux inmux_16_13_65813_65823 (
    .I(net_65813),
    .O(net_65823)
  );
  InMux inmux_16_13_65814_65853 (
    .I(net_65814),
    .O(net_65853)
  );
  InMux inmux_16_13_65815_65866 (
    .I(net_65815),
    .O(net_65866)
  );
  InMux inmux_16_13_65816_65841 (
    .I(net_65816),
    .O(net_65841)
  );
  InMux inmux_16_13_65819_65852 (
    .I(net_65819),
    .O(net_65852)
  );
  InMux inmux_16_13_65820_65830 (
    .I(net_65820),
    .O(net_65830)
  );
  InMux inmux_16_13_65826_65836 (
    .I(net_65826),
    .O(net_65836)
  );
  InMux inmux_16_13_65832_65842 (
    .I(net_65832),
    .O(net_65842)
  );
  InMux inmux_16_13_65838_65848 (
    .I(net_65838),
    .O(net_65848)
  );
  InMux inmux_16_13_65844_65854 (
    .I(net_65844),
    .O(net_65854)
  );
  InMux inmux_16_13_65850_65860 (
    .I(net_65850),
    .O(net_65860)
  );
  SRMux inmux_16_13_9_65869 (
    .I(net_9),
    .O(net_65869)
  );
  InMux inmux_16_14_65911_65963 (
    .I(net_65911),
    .O(net_65963)
  );
  InMux inmux_16_14_65912_65952 (
    .I(net_65912),
    .O(net_65952)
  );
  InMux inmux_16_14_65913_65975 (
    .I(net_65913),
    .O(net_65975)
  );
  InMux inmux_16_14_65917_65987 (
    .I(net_65917),
    .O(net_65987)
  );
  InMux inmux_16_14_65919_65976 (
    .I(net_65919),
    .O(net_65976)
  );
  InMux inmux_16_14_65923_65981 (
    .I(net_65923),
    .O(net_65981)
  );
  InMux inmux_16_14_65924_65982 (
    .I(net_65924),
    .O(net_65982)
  );
  InMux inmux_16_14_65925_65969 (
    .I(net_65925),
    .O(net_65969)
  );
  InMux inmux_16_14_65926_65958 (
    .I(net_65926),
    .O(net_65958)
  );
  InMux inmux_16_14_65930_65964 (
    .I(net_65930),
    .O(net_65964)
  );
  InMux inmux_16_14_65933_65951 (
    .I(net_65933),
    .O(net_65951)
  );
  InMux inmux_16_14_65934_65945 (
    .I(net_65934),
    .O(net_65945)
  );
  InMux inmux_16_14_65935_65988 (
    .I(net_65935),
    .O(net_65988)
  );
  InMux inmux_16_14_65937_65957 (
    .I(net_65937),
    .O(net_65957)
  );
  InMux inmux_16_14_65938_65970 (
    .I(net_65938),
    .O(net_65970)
  );
  InMux inmux_16_14_65940_65946 (
    .I(net_65940),
    .O(net_65946)
  );
  InMux inmux_16_14_65943_65953 (
    .I(net_65943),
    .O(net_65953)
  );
  InMux inmux_16_14_65949_65959 (
    .I(net_65949),
    .O(net_65959)
  );
  InMux inmux_16_14_65955_65965 (
    .I(net_65955),
    .O(net_65965)
  );
  InMux inmux_16_14_65961_65971 (
    .I(net_65961),
    .O(net_65971)
  );
  InMux inmux_16_14_65967_65977 (
    .I(net_65967),
    .O(net_65977)
  );
  InMux inmux_16_14_65973_65983 (
    .I(net_65973),
    .O(net_65983)
  );
  InMux inmux_16_14_65979_65989 (
    .I(net_65979),
    .O(net_65989)
  );
  ClkMux inmux_16_15_5_66114 (
    .I(net_5),
    .O(net_66114)
  );
  InMux inmux_16_15_66029_66070 (
    .I(net_66029),
    .O(net_66070)
  );
  InMux inmux_16_15_66040_66067 (
    .I(net_66040),
    .O(net_66067)
  );
  InMux inmux_16_15_66041_66092 (
    .I(net_66041),
    .O(net_66092)
  );
  InMux inmux_16_15_66049_66100 (
    .I(net_66049),
    .O(net_66100)
  );
  InMux inmux_16_15_66050_66105 (
    .I(net_66050),
    .O(net_66105)
  );
  InMux inmux_16_15_66051_66075 (
    .I(net_66051),
    .O(net_66075)
  );
  InMux inmux_16_15_66054_66069 (
    .I(net_66054),
    .O(net_66069)
  );
  InMux inmux_16_15_66063_66086 (
    .I(net_66063),
    .O(net_66086)
  );
  InMux inmux_16_15_66063_66112 (
    .I(net_66063),
    .O(net_66112)
  );
  InMux inmux_16_15_66064_66080 (
    .I(net_66064),
    .O(net_66080)
  );
  SRMux inmux_16_15_9_66115 (
    .I(net_9),
    .O(net_66115)
  );
  ClkMux inmux_16_16_5_66237 (
    .I(net_5),
    .O(net_66237)
  );
  InMux inmux_16_16_66160_66191 (
    .I(net_66160),
    .O(net_66191)
  );
  InMux inmux_16_16_66161_66223 (
    .I(net_66161),
    .O(net_66223)
  );
  InMux inmux_16_16_66162_66227 (
    .I(net_66162),
    .O(net_66227)
  );
  InMux inmux_16_16_66164_66205 (
    .I(net_66164),
    .O(net_66205)
  );
  InMux inmux_16_16_66165_66210 (
    .I(net_66165),
    .O(net_66210)
  );
  InMux inmux_16_16_66167_66198 (
    .I(net_66167),
    .O(net_66198)
  );
  InMux inmux_16_16_66169_66193 (
    .I(net_66169),
    .O(net_66193)
  );
  InMux inmux_16_16_66171_66229 (
    .I(net_66171),
    .O(net_66229)
  );
  InMux inmux_16_16_66172_66190 (
    .I(net_66172),
    .O(net_66190)
  );
  InMux inmux_16_16_66172_66199 (
    .I(net_66172),
    .O(net_66199)
  );
  InMux inmux_16_16_66172_66202 (
    .I(net_66172),
    .O(net_66202)
  );
  InMux inmux_16_16_66172_66228 (
    .I(net_66172),
    .O(net_66228)
  );
  InMux inmux_16_16_66176_66234 (
    .I(net_66176),
    .O(net_66234)
  );
  InMux inmux_16_16_66180_66215 (
    .I(net_66180),
    .O(net_66215)
  );
  InMux inmux_16_16_66185_66196 (
    .I(net_66185),
    .O(net_66196)
  );
  InMux inmux_16_16_66187_66203 (
    .I(net_66187),
    .O(net_66203)
  );
  InMux inmux_16_16_66188_66192 (
    .I(net_66188),
    .O(net_66192)
  );
  InMux inmux_16_16_66188_66197 (
    .I(net_66188),
    .O(net_66197)
  );
  InMux inmux_16_16_66188_66204 (
    .I(net_66188),
    .O(net_66204)
  );
  InMux inmux_16_16_66188_66209 (
    .I(net_66188),
    .O(net_66209)
  );
  InMux inmux_16_16_66188_66216 (
    .I(net_66188),
    .O(net_66216)
  );
  InMux inmux_16_16_66188_66221 (
    .I(net_66188),
    .O(net_66221)
  );
  InMux inmux_16_16_66188_66226 (
    .I(net_66188),
    .O(net_66226)
  );
  InMux inmux_16_16_66188_66235 (
    .I(net_66188),
    .O(net_66235)
  );
  CEMux inmux_16_16_6_66236 (
    .I(net_6),
    .O(net_66236)
  );
  SRMux inmux_16_16_9_66238 (
    .I(net_9),
    .O(net_66238)
  );
  ClkMux inmux_16_17_5_66360 (
    .I(net_5),
    .O(net_66360)
  );
  InMux inmux_16_17_66280_66356 (
    .I(net_66280),
    .O(net_66356)
  );
  InMux inmux_16_17_66282_66332 (
    .I(net_66282),
    .O(net_66332)
  );
  InMux inmux_16_17_66283_66331 (
    .I(net_66283),
    .O(net_66331)
  );
  InMux inmux_16_17_66284_66327 (
    .I(net_66284),
    .O(net_66327)
  );
  InMux inmux_16_17_66293_66315 (
    .I(net_66293),
    .O(net_66315)
  );
  InMux inmux_16_17_66297_66326 (
    .I(net_66297),
    .O(net_66326)
  );
  InMux inmux_16_17_66299_66321 (
    .I(net_66299),
    .O(net_66321)
  );
  InMux inmux_16_17_66302_66325 (
    .I(net_66302),
    .O(net_66325)
  );
  InMux inmux_16_17_66302_66358 (
    .I(net_66302),
    .O(net_66358)
  );
  InMux inmux_16_17_66303_66314 (
    .I(net_66303),
    .O(net_66314)
  );
  InMux inmux_16_17_66303_66319 (
    .I(net_66303),
    .O(net_66319)
  );
  InMux inmux_16_17_66303_66328 (
    .I(net_66303),
    .O(net_66328)
  );
  InMux inmux_16_17_66303_66338 (
    .I(net_66303),
    .O(net_66338)
  );
  InMux inmux_16_17_66303_66345 (
    .I(net_66303),
    .O(net_66345)
  );
  InMux inmux_16_17_66303_66350 (
    .I(net_66303),
    .O(net_66350)
  );
  InMux inmux_16_17_66303_66357 (
    .I(net_66303),
    .O(net_66357)
  );
  InMux inmux_16_17_66304_66355 (
    .I(net_66304),
    .O(net_66355)
  );
  InMux inmux_16_17_66305_66349 (
    .I(net_66305),
    .O(net_66349)
  );
  InMux inmux_16_17_66308_66343 (
    .I(net_66308),
    .O(net_66343)
  );
  InMux inmux_16_17_66310_66340 (
    .I(net_66310),
    .O(net_66340)
  );
  CEMux inmux_16_17_6_66359 (
    .I(net_6),
    .O(net_66359)
  );
  SRMux inmux_16_17_9_66361 (
    .I(net_9),
    .O(net_66361)
  );
  ClkMux inmux_16_18_5_66483 (
    .I(net_5),
    .O(net_66483)
  );
  CEMux inmux_16_18_66414_66482 (
    .I(net_66414),
    .O(net_66482)
  );
  InMux inmux_16_18_66425_66438 (
    .I(net_66425),
    .O(net_66438)
  );
  SRMux inmux_16_18_9_66484 (
    .I(net_9),
    .O(net_66484)
  );
  CEMux inmux_16_2_10_64514 (
    .I(net_10),
    .O(net_64514)
  );
  ClkMux inmux_16_2_5_64515 (
    .I(net_5),
    .O(net_64515)
  );
  InMux inmux_16_2_64440_64488 (
    .I(net_64440),
    .O(net_64488)
  );
  IoInMux inmux_16_31_68021_68006 (
    .I(net_68021),
    .O(net_68006)
  );
  IoInMux inmux_16_31_68025_68009 (
    .I(net_68025),
    .O(net_68009)
  );
  ClkMux inmux_16_3_5_64638 (
    .I(net_5),
    .O(net_64638)
  );
  CEMux inmux_16_3_64560_64637 (
    .I(net_64560),
    .O(net_64637)
  );
  InMux inmux_16_3_64564_64610 (
    .I(net_64564),
    .O(net_64610)
  );
  InMux inmux_16_3_64568_64604 (
    .I(net_64568),
    .O(net_64604)
  );
  InMux inmux_16_3_64569_64603 (
    .I(net_64569),
    .O(net_64603)
  );
  InMux inmux_16_3_64580_64605 (
    .I(net_64580),
    .O(net_64605)
  );
  InMux inmux_16_3_64585_64612 (
    .I(net_64585),
    .O(net_64612)
  );
  InMux inmux_16_3_64586_64606 (
    .I(net_64586),
    .O(net_64606)
  );
  SRMux inmux_16_3_9_64639 (
    .I(net_9),
    .O(net_64639)
  );
  InMux inmux_16_4_64685_64728 (
    .I(net_64685),
    .O(net_64728)
  );
  InMux inmux_16_4_64688_64758 (
    .I(net_64688),
    .O(net_64758)
  );
  InMux inmux_16_4_64692_64721 (
    .I(net_64692),
    .O(net_64721)
  );
  InMux inmux_16_4_64693_64746 (
    .I(net_64693),
    .O(net_64746)
  );
  InMux inmux_16_4_64695_64734 (
    .I(net_64695),
    .O(net_64734)
  );
  InMux inmux_16_4_64696_64757 (
    .I(net_64696),
    .O(net_64757)
  );
  InMux inmux_16_4_64697_64716 (
    .I(net_64697),
    .O(net_64716)
  );
  InMux inmux_16_4_64698_64727 (
    .I(net_64698),
    .O(net_64727)
  );
  InMux inmux_16_4_64699_64752 (
    .I(net_64699),
    .O(net_64752)
  );
  InMux inmux_16_4_64700_64739 (
    .I(net_64700),
    .O(net_64739)
  );
  InMux inmux_16_4_64701_64745 (
    .I(net_64701),
    .O(net_64745)
  );
  InMux inmux_16_4_64702_64722 (
    .I(net_64702),
    .O(net_64722)
  );
  InMux inmux_16_4_64703_64740 (
    .I(net_64703),
    .O(net_64740)
  );
  InMux inmux_16_4_64705_64751 (
    .I(net_64705),
    .O(net_64751)
  );
  InMux inmux_16_4_64711_64715 (
    .I(net_64711),
    .O(net_64715)
  );
  InMux inmux_16_4_64712_64733 (
    .I(net_64712),
    .O(net_64733)
  );
  InMux inmux_16_4_64713_64723 (
    .I(net_64713),
    .O(net_64723)
  );
  InMux inmux_16_4_64719_64729 (
    .I(net_64719),
    .O(net_64729)
  );
  InMux inmux_16_4_64725_64735 (
    .I(net_64725),
    .O(net_64735)
  );
  InMux inmux_16_4_64731_64741 (
    .I(net_64731),
    .O(net_64741)
  );
  InMux inmux_16_4_64737_64747 (
    .I(net_64737),
    .O(net_64747)
  );
  InMux inmux_16_4_64743_64753 (
    .I(net_64743),
    .O(net_64753)
  );
  InMux inmux_16_4_64749_64759 (
    .I(net_64749),
    .O(net_64759)
  );
  ClkMux inmux_16_5_5_64884 (
    .I(net_5),
    .O(net_64884)
  );
  InMux inmux_16_5_64799_64840 (
    .I(net_64799),
    .O(net_64840)
  );
  InMux inmux_16_5_64805_64881 (
    .I(net_64805),
    .O(net_64881)
  );
  InMux inmux_16_5_64812_64876 (
    .I(net_64812),
    .O(net_64876)
  );
  InMux inmux_16_5_64817_64861 (
    .I(net_64817),
    .O(net_64861)
  );
  InMux inmux_16_5_64820_64868 (
    .I(net_64820),
    .O(net_64868)
  );
  InMux inmux_16_5_64822_64851 (
    .I(net_64822),
    .O(net_64851)
  );
  InMux inmux_16_5_64823_64850 (
    .I(net_64823),
    .O(net_64850)
  );
  InMux inmux_16_5_64826_64870 (
    .I(net_64826),
    .O(net_64870)
  );
  InMux inmux_16_5_64829_64839 (
    .I(net_64829),
    .O(net_64839)
  );
  InMux inmux_16_5_64830_64845 (
    .I(net_64830),
    .O(net_64845)
  );
  InMux inmux_16_5_64834_64838 (
    .I(net_64834),
    .O(net_64838)
  );
  InMux inmux_16_5_64835_64844 (
    .I(net_64835),
    .O(net_64844)
  );
  InMux inmux_16_5_64836_64846 (
    .I(net_64836),
    .O(net_64846)
  );
  InMux inmux_16_5_64842_64852 (
    .I(net_64842),
    .O(net_64852)
  );
  InMux inmux_16_5_64848_64858 (
    .I(net_64848),
    .O(net_64858)
  );
  SRMux inmux_16_5_9_64885 (
    .I(net_9),
    .O(net_64885)
  );
  ClkMux inmux_16_6_5_65007 (
    .I(net_5),
    .O(net_65007)
  );
  InMux inmux_16_6_64929_64962 (
    .I(net_64929),
    .O(net_64962)
  );
  InMux inmux_16_6_64931_64974 (
    .I(net_64931),
    .O(net_64974)
  );
  InMux inmux_16_6_64932_64961 (
    .I(net_64932),
    .O(net_64961)
  );
  InMux inmux_16_6_64933_64979 (
    .I(net_64933),
    .O(net_64979)
  );
  InMux inmux_16_6_64938_64991 (
    .I(net_64938),
    .O(net_64991)
  );
  InMux inmux_16_6_64941_65004 (
    .I(net_64941),
    .O(net_65004)
  );
  InMux inmux_16_6_64946_64968 (
    .I(net_64946),
    .O(net_64968)
  );
  InMux inmux_16_6_64952_64986 (
    .I(net_64952),
    .O(net_64986)
  );
  InMux inmux_16_6_64956_64998 (
    .I(net_64956),
    .O(net_64998)
  );
  InMux inmux_16_6_64959_64969 (
    .I(net_64959),
    .O(net_64969)
  );
  InMux inmux_16_6_64965_64975 (
    .I(net_64965),
    .O(net_64975)
  );
  InMux inmux_16_6_64971_64981 (
    .I(net_64971),
    .O(net_64981)
  );
  InMux inmux_16_6_64977_64987 (
    .I(net_64977),
    .O(net_64987)
  );
  InMux inmux_16_6_64983_64993 (
    .I(net_64983),
    .O(net_64993)
  );
  InMux inmux_16_6_64989_64999 (
    .I(net_64989),
    .O(net_64999)
  );
  InMux inmux_16_6_64995_65005 (
    .I(net_64995),
    .O(net_65005)
  );
  SRMux inmux_16_6_9_65008 (
    .I(net_9),
    .O(net_65008)
  );
  ClkMux inmux_16_7_5_65130 (
    .I(net_5),
    .O(net_65130)
  );
  InMux inmux_16_7_65045_65086 (
    .I(net_65045),
    .O(net_65086)
  );
  InMux inmux_16_7_65050_65085 (
    .I(net_65050),
    .O(net_65085)
  );
  InMux inmux_16_7_65052_65090 (
    .I(net_65052),
    .O(net_65090)
  );
  InMux inmux_16_7_65053_65122 (
    .I(net_65053),
    .O(net_65122)
  );
  InMux inmux_16_7_65054_65116 (
    .I(net_65054),
    .O(net_65116)
  );
  InMux inmux_16_7_65062_65096 (
    .I(net_65062),
    .O(net_65096)
  );
  InMux inmux_16_7_65065_65121 (
    .I(net_65065),
    .O(net_65121)
  );
  InMux inmux_16_7_65070_65126 (
    .I(net_65070),
    .O(net_65126)
  );
  InMux inmux_16_7_65073_65103 (
    .I(net_65073),
    .O(net_65103)
  );
  InMux inmux_16_7_65082_65092 (
    .I(net_65082),
    .O(net_65092)
  );
  InMux inmux_16_7_65088_65098 (
    .I(net_65088),
    .O(net_65098)
  );
  InMux inmux_16_7_65094_65104 (
    .I(net_65094),
    .O(net_65104)
  );
  InMux inmux_16_7_65100_65110 (
    .I(net_65100),
    .O(net_65110)
  );
  SRMux inmux_16_7_9_65131 (
    .I(net_9),
    .O(net_65131)
  );
  ClkMux inmux_16_8_5_65253 (
    .I(net_5),
    .O(net_65253)
  );
  InMux inmux_16_8_65176_65207 (
    .I(net_65176),
    .O(net_65207)
  );
  InMux inmux_16_8_65180_65214 (
    .I(net_65180),
    .O(net_65214)
  );
  InMux inmux_16_8_65185_65212 (
    .I(net_65185),
    .O(net_65212)
  );
  InMux inmux_16_8_65186_65232 (
    .I(net_65186),
    .O(net_65232)
  );
  SRMux inmux_16_8_9_65254 (
    .I(net_9),
    .O(net_65254)
  );
  ClkMux inmux_16_9_5_65376 (
    .I(net_5),
    .O(net_65376)
  );
  InMux inmux_16_9_65303_65337 (
    .I(net_65303),
    .O(net_65337)
  );
  InMux inmux_16_9_65304_65356 (
    .I(net_65304),
    .O(net_65356)
  );
  InMux inmux_16_9_65307_65362 (
    .I(net_65307),
    .O(net_65362)
  );
  InMux inmux_16_9_65310_65366 (
    .I(net_65310),
    .O(net_65366)
  );
  InMux inmux_16_9_65319_65344 (
    .I(net_65319),
    .O(net_65344)
  );
  InMux inmux_16_9_65327_65372 (
    .I(net_65327),
    .O(net_65372)
  );
  SRMux inmux_16_9_9_65377 (
    .I(net_9),
    .O(net_65377)
  );
  ClkMux inmux_17_10_5_69330 (
    .I(net_5),
    .O(net_69330)
  );
  InMux inmux_17_10_69254_69295 (
    .I(net_69254),
    .O(net_69295)
  );
  InMux inmux_17_10_69258_69303 (
    .I(net_69258),
    .O(net_69303)
  );
  InMux inmux_17_10_69263_69316 (
    .I(net_69263),
    .O(net_69316)
  );
  InMux inmux_17_10_69265_69292 (
    .I(net_69265),
    .O(net_69292)
  );
  InMux inmux_17_10_69269_69286 (
    .I(net_69269),
    .O(net_69286)
  );
  InMux inmux_17_10_69270_69326 (
    .I(net_69270),
    .O(net_69326)
  );
  InMux inmux_17_10_69280_69308 (
    .I(net_69280),
    .O(net_69308)
  );
  SRMux inmux_17_10_9_69331 (
    .I(net_9),
    .O(net_69331)
  );
  ClkMux inmux_17_11_5_69453 (
    .I(net_5),
    .O(net_69453)
  );
  InMux inmux_17_11_69373_69449 (
    .I(net_69373),
    .O(net_69449)
  );
  InMux inmux_17_11_69374_69407 (
    .I(net_69374),
    .O(net_69407)
  );
  InMux inmux_17_11_69378_69438 (
    .I(net_69378),
    .O(net_69438)
  );
  InMux inmux_17_11_69380_69445 (
    .I(net_69380),
    .O(net_69445)
  );
  InMux inmux_17_11_69380_69448 (
    .I(net_69380),
    .O(net_69448)
  );
  InMux inmux_17_11_69381_69414 (
    .I(net_69381),
    .O(net_69414)
  );
  CEMux inmux_17_11_69384_69452 (
    .I(net_69384),
    .O(net_69452)
  );
  InMux inmux_17_11_69385_69426 (
    .I(net_69385),
    .O(net_69426)
  );
  InMux inmux_17_11_69386_69437 (
    .I(net_69386),
    .O(net_69437)
  );
  InMux inmux_17_11_69388_69413 (
    .I(net_69388),
    .O(net_69413)
  );
  InMux inmux_17_11_69389_69420 (
    .I(net_69389),
    .O(net_69420)
  );
  InMux inmux_17_11_69391_69425 (
    .I(net_69391),
    .O(net_69425)
  );
  InMux inmux_17_11_69395_69408 (
    .I(net_69395),
    .O(net_69408)
  );
  InMux inmux_17_11_69397_69431 (
    .I(net_69397),
    .O(net_69431)
  );
  InMux inmux_17_11_69399_69436 (
    .I(net_69399),
    .O(net_69436)
  );
  InMux inmux_17_11_69402_69442 (
    .I(net_69402),
    .O(net_69442)
  );
  InMux inmux_17_11_69403_69419 (
    .I(net_69403),
    .O(net_69419)
  );
  InMux inmux_17_11_69405_69415 (
    .I(net_69405),
    .O(net_69415)
  );
  InMux inmux_17_11_69411_69421 (
    .I(net_69411),
    .O(net_69421)
  );
  InMux inmux_17_11_69417_69427 (
    .I(net_69417),
    .O(net_69427)
  );
  InMux inmux_17_11_69423_69433 (
    .I(net_69423),
    .O(net_69433)
  );
  InMux inmux_17_11_69429_69439 (
    .I(net_69429),
    .O(net_69439)
  );
  SRMux inmux_17_11_9_69454 (
    .I(net_9),
    .O(net_69454)
  );
  ClkMux inmux_17_12_5_69576 (
    .I(net_5),
    .O(net_69576)
  );
  InMux inmux_17_12_69499_69532 (
    .I(net_69499),
    .O(net_69532)
  );
  InMux inmux_17_12_69509_69560 (
    .I(net_69509),
    .O(net_69560)
  );
  InMux inmux_17_12_69515_69535 (
    .I(net_69515),
    .O(net_69535)
  );
  InMux inmux_17_12_69518_69574 (
    .I(net_69518),
    .O(net_69574)
  );
  InMux inmux_17_12_69521_69541 (
    .I(net_69521),
    .O(net_69541)
  );
  InMux inmux_17_12_69522_69549 (
    .I(net_69522),
    .O(net_69549)
  );
  InMux inmux_17_12_69525_69555 (
    .I(net_69525),
    .O(net_69555)
  );
  InMux inmux_17_12_69526_69568 (
    .I(net_69526),
    .O(net_69568)
  );
  SRMux inmux_17_12_9_69577 (
    .I(net_9),
    .O(net_69577)
  );
  InMux inmux_17_13_69623_69654 (
    .I(net_69623),
    .O(net_69654)
  );
  InMux inmux_17_13_69637_69666 (
    .I(net_69637),
    .O(net_69666)
  );
  InMux inmux_17_13_69638_69653 (
    .I(net_69638),
    .O(net_69653)
  );
  InMux inmux_17_13_69638_69660 (
    .I(net_69638),
    .O(net_69660)
  );
  InMux inmux_17_13_69638_69665 (
    .I(net_69638),
    .O(net_69665)
  );
  InMux inmux_17_13_69638_69672 (
    .I(net_69638),
    .O(net_69672)
  );
  InMux inmux_17_13_69638_69677 (
    .I(net_69638),
    .O(net_69677)
  );
  InMux inmux_17_13_69638_69684 (
    .I(net_69638),
    .O(net_69684)
  );
  InMux inmux_17_13_69638_69689 (
    .I(net_69638),
    .O(net_69689)
  );
  InMux inmux_17_13_69638_69696 (
    .I(net_69638),
    .O(net_69696)
  );
  InMux inmux_17_13_69639_69678 (
    .I(net_69639),
    .O(net_69678)
  );
  InMux inmux_17_13_69641_69690 (
    .I(net_69641),
    .O(net_69690)
  );
  InMux inmux_17_13_69644_69659 (
    .I(net_69644),
    .O(net_69659)
  );
  InMux inmux_17_13_69646_69671 (
    .I(net_69646),
    .O(net_69671)
  );
  InMux inmux_17_13_69648_69683 (
    .I(net_69648),
    .O(net_69683)
  );
  InMux inmux_17_13_69650_69695 (
    .I(net_69650),
    .O(net_69695)
  );
  InMux inmux_17_13_69651_69661 (
    .I(net_69651),
    .O(net_69661)
  );
  InMux inmux_17_13_69657_69667 (
    .I(net_69657),
    .O(net_69667)
  );
  InMux inmux_17_13_69663_69673 (
    .I(net_69663),
    .O(net_69673)
  );
  InMux inmux_17_13_69669_69679 (
    .I(net_69669),
    .O(net_69679)
  );
  InMux inmux_17_13_69675_69685 (
    .I(net_69675),
    .O(net_69685)
  );
  InMux inmux_17_13_69681_69691 (
    .I(net_69681),
    .O(net_69691)
  );
  ClkMux inmux_17_14_5_69822 (
    .I(net_5),
    .O(net_69822)
  );
  InMux inmux_17_14_69737_69778 (
    .I(net_69737),
    .O(net_69778)
  );
  InMux inmux_17_14_69744_69794 (
    .I(net_69744),
    .O(net_69794)
  );
  InMux inmux_17_14_69746_69808 (
    .I(net_69746),
    .O(net_69808)
  );
  InMux inmux_17_14_69747_69788 (
    .I(net_69747),
    .O(net_69788)
  );
  InMux inmux_17_14_69747_69795 (
    .I(net_69747),
    .O(net_69795)
  );
  InMux inmux_17_14_69747_69812 (
    .I(net_69747),
    .O(net_69812)
  );
  InMux inmux_17_14_69748_69784 (
    .I(net_69748),
    .O(net_69784)
  );
  InMux inmux_17_14_69748_69818 (
    .I(net_69748),
    .O(net_69818)
  );
  InMux inmux_17_14_69753_69813 (
    .I(net_69753),
    .O(net_69813)
  );
  InMux inmux_17_14_69754_69781 (
    .I(net_69754),
    .O(net_69781)
  );
  InMux inmux_17_14_69755_69787 (
    .I(net_69755),
    .O(net_69787)
  );
  InMux inmux_17_14_69756_69817 (
    .I(net_69756),
    .O(net_69817)
  );
  InMux inmux_17_14_69757_69799 (
    .I(net_69757),
    .O(net_69799)
  );
  InMux inmux_17_14_69758_69775 (
    .I(net_69758),
    .O(net_69775)
  );
  InMux inmux_17_14_69760_69801 (
    .I(net_69760),
    .O(net_69801)
  );
  InMux inmux_17_14_69762_69796 (
    .I(net_69762),
    .O(net_69796)
  );
  InMux inmux_17_14_69763_69800 (
    .I(net_69763),
    .O(net_69800)
  );
  InMux inmux_17_14_69764_69777 (
    .I(net_69764),
    .O(net_69777)
  );
  InMux inmux_17_14_69765_69793 (
    .I(net_69765),
    .O(net_69793)
  );
  InMux inmux_17_14_69766_69783 (
    .I(net_69766),
    .O(net_69783)
  );
  InMux inmux_17_14_69768_69790 (
    .I(net_69768),
    .O(net_69790)
  );
  InMux inmux_17_14_69770_69819 (
    .I(net_69770),
    .O(net_69819)
  );
  InMux inmux_17_14_69772_69814 (
    .I(net_69772),
    .O(net_69814)
  );
  InMux inmux_17_14_69773_69782 (
    .I(net_69773),
    .O(net_69782)
  );
  InMux inmux_17_14_69773_69789 (
    .I(net_69773),
    .O(net_69789)
  );
  InMux inmux_17_14_69773_69811 (
    .I(net_69773),
    .O(net_69811)
  );
  InMux inmux_17_14_69773_69820 (
    .I(net_69773),
    .O(net_69820)
  );
  CEMux inmux_17_14_6_69821 (
    .I(net_6),
    .O(net_69821)
  );
  SRMux inmux_17_14_9_69823 (
    .I(net_9),
    .O(net_69823)
  );
  ClkMux inmux_17_15_5_69945 (
    .I(net_5),
    .O(net_69945)
  );
  InMux inmux_17_15_69868_69911 (
    .I(net_69868),
    .O(net_69911)
  );
  InMux inmux_17_15_69882_69930 (
    .I(net_69882),
    .O(net_69930)
  );
  InMux inmux_17_15_69883_69900 (
    .I(net_69883),
    .O(net_69900)
  );
  InMux inmux_17_15_69884_69925 (
    .I(net_69884),
    .O(net_69925)
  );
  InMux inmux_17_15_69886_69918 (
    .I(net_69886),
    .O(net_69918)
  );
  InMux inmux_17_15_69891_69940 (
    .I(net_69891),
    .O(net_69940)
  );
  InMux inmux_17_15_69892_69934 (
    .I(net_69892),
    .O(net_69934)
  );
  InMux inmux_17_15_69894_69905 (
    .I(net_69894),
    .O(net_69905)
  );
  SRMux inmux_17_15_9_69946 (
    .I(net_9),
    .O(net_69946)
  );
  InMux inmux_17_16_69990_70035 (
    .I(net_69990),
    .O(net_70035)
  );
  InMux inmux_17_16_69991_70041 (
    .I(net_69991),
    .O(net_70041)
  );
  InMux inmux_17_16_69997_70028 (
    .I(net_69997),
    .O(net_70028)
  );
  InMux inmux_17_16_70000_70046 (
    .I(net_70000),
    .O(net_70046)
  );
  InMux inmux_17_16_70001_70052 (
    .I(net_70001),
    .O(net_70052)
  );
  InMux inmux_17_16_70002_70058 (
    .I(net_70002),
    .O(net_70058)
  );
  InMux inmux_17_16_70003_70064 (
    .I(net_70003),
    .O(net_70064)
  );
  InMux inmux_17_16_70008_70023 (
    .I(net_70008),
    .O(net_70023)
  );
  InMux inmux_17_16_70016_70022 (
    .I(net_70016),
    .O(net_70022)
  );
  InMux inmux_17_16_70020_70030 (
    .I(net_70020),
    .O(net_70030)
  );
  InMux inmux_17_16_70026_70036 (
    .I(net_70026),
    .O(net_70036)
  );
  InMux inmux_17_16_70032_70042 (
    .I(net_70032),
    .O(net_70042)
  );
  InMux inmux_17_16_70038_70048 (
    .I(net_70038),
    .O(net_70048)
  );
  InMux inmux_17_16_70044_70054 (
    .I(net_70044),
    .O(net_70054)
  );
  InMux inmux_17_16_70050_70060 (
    .I(net_70050),
    .O(net_70060)
  );
  ClkMux inmux_17_17_5_70191 (
    .I(net_5),
    .O(net_70191)
  );
  CEMux inmux_17_17_6_70190 (
    .I(net_6),
    .O(net_70190)
  );
  InMux inmux_17_17_70106_70147 (
    .I(net_70106),
    .O(net_70147)
  );
  InMux inmux_17_17_70111_70168 (
    .I(net_70111),
    .O(net_70168)
  );
  InMux inmux_17_17_70111_70187 (
    .I(net_70111),
    .O(net_70187)
  );
  InMux inmux_17_17_70114_70169 (
    .I(net_70114),
    .O(net_70169)
  );
  InMux inmux_17_17_70114_70186 (
    .I(net_70114),
    .O(net_70186)
  );
  InMux inmux_17_17_70115_70163 (
    .I(net_70115),
    .O(net_70163)
  );
  InMux inmux_17_17_70116_70152 (
    .I(net_70116),
    .O(net_70152)
  );
  InMux inmux_17_17_70117_70151 (
    .I(net_70117),
    .O(net_70151)
  );
  InMux inmux_17_17_70117_70170 (
    .I(net_70117),
    .O(net_70170)
  );
  InMux inmux_17_17_70117_70182 (
    .I(net_70117),
    .O(net_70182)
  );
  InMux inmux_17_17_70117_70189 (
    .I(net_70117),
    .O(net_70189)
  );
  InMux inmux_17_17_70118_70150 (
    .I(net_70118),
    .O(net_70150)
  );
  InMux inmux_17_17_70118_70171 (
    .I(net_70118),
    .O(net_70171)
  );
  InMux inmux_17_17_70118_70181 (
    .I(net_70118),
    .O(net_70181)
  );
  InMux inmux_17_17_70118_70188 (
    .I(net_70118),
    .O(net_70188)
  );
  InMux inmux_17_17_70119_70183 (
    .I(net_70119),
    .O(net_70183)
  );
  InMux inmux_17_17_70120_70180 (
    .I(net_70120),
    .O(net_70180)
  );
  InMux inmux_17_17_70124_70177 (
    .I(net_70124),
    .O(net_70177)
  );
  InMux inmux_17_17_70131_70165 (
    .I(net_70131),
    .O(net_70165)
  );
  InMux inmux_17_17_70134_70174 (
    .I(net_70134),
    .O(net_70174)
  );
  InMux inmux_17_17_70138_70153 (
    .I(net_70138),
    .O(net_70153)
  );
  SRMux inmux_17_17_9_70192 (
    .I(net_9),
    .O(net_70192)
  );
  ClkMux inmux_17_18_5_70314 (
    .I(net_5),
    .O(net_70314)
  );
  InMux inmux_17_18_70238_70303 (
    .I(net_70238),
    .O(net_70303)
  );
  SRMux inmux_17_18_9_70315 (
    .I(net_9),
    .O(net_70315)
  );
  CEMux inmux_17_2_10_68345 (
    .I(net_10),
    .O(net_68345)
  );
  ClkMux inmux_17_2_5_68346 (
    .I(net_5),
    .O(net_68346)
  );
  InMux inmux_17_2_68281_68299 (
    .I(net_68281),
    .O(net_68299)
  );
  InMux inmux_17_2_68292_68341 (
    .I(net_68292),
    .O(net_68341)
  );
  IoInMux inmux_17_31_71855_71837 (
    .I(net_71855),
    .O(net_71837)
  );
  ClkMux inmux_17_3_5_68469 (
    .I(net_5),
    .O(net_68469)
  );
  InMux inmux_17_3_68391_68436 (
    .I(net_68391),
    .O(net_68436)
  );
  InMux inmux_17_3_68392_68430 (
    .I(net_68392),
    .O(net_68430)
  );
  InMux inmux_17_3_68400_68446 (
    .I(net_68400),
    .O(net_68446)
  );
  InMux inmux_17_3_68409_68424 (
    .I(net_68409),
    .O(net_68424)
  );
  InMux inmux_17_3_68413_68440 (
    .I(net_68413),
    .O(net_68440)
  );
  SRMux inmux_17_3_9_68470 (
    .I(net_9),
    .O(net_68470)
  );
  ClkMux inmux_17_4_5_68592 (
    .I(net_5),
    .O(net_68592)
  );
  InMux inmux_17_4_68515_68560 (
    .I(net_68515),
    .O(net_68560)
  );
  InMux inmux_17_4_68520_68589 (
    .I(net_68520),
    .O(net_68589)
  );
  InMux inmux_17_4_68522_68553 (
    .I(net_68522),
    .O(net_68553)
  );
  InMux inmux_17_4_68523_68583 (
    .I(net_68523),
    .O(net_68583)
  );
  InMux inmux_17_4_68525_68578 (
    .I(net_68525),
    .O(net_68578)
  );
  InMux inmux_17_4_68526_68572 (
    .I(net_68526),
    .O(net_68572)
  );
  InMux inmux_17_4_68527_68566 (
    .I(net_68527),
    .O(net_68566)
  );
  InMux inmux_17_4_68535_68546 (
    .I(net_68535),
    .O(net_68546)
  );
  SRMux inmux_17_4_9_68593 (
    .I(net_9),
    .O(net_68593)
  );
  ClkMux inmux_17_5_5_68715 (
    .I(net_5),
    .O(net_68715)
  );
  InMux inmux_17_5_68638_68674 (
    .I(net_68638),
    .O(net_68674)
  );
  InMux inmux_17_5_68642_68698 (
    .I(net_68642),
    .O(net_68698)
  );
  InMux inmux_17_5_68643_68712 (
    .I(net_68643),
    .O(net_68712)
  );
  InMux inmux_17_5_68644_68706 (
    .I(net_68644),
    .O(net_68706)
  );
  InMux inmux_17_5_68646_68687 (
    .I(net_68646),
    .O(net_68687)
  );
  InMux inmux_17_5_68653_68682 (
    .I(net_68653),
    .O(net_68682)
  );
  InMux inmux_17_5_68666_68670 (
    .I(net_68666),
    .O(net_68670)
  );
  SRMux inmux_17_5_9_68716 (
    .I(net_9),
    .O(net_68716)
  );
  ClkMux inmux_17_6_5_68838 (
    .I(net_5),
    .O(net_68838)
  );
  InMux inmux_17_6_68764_68805 (
    .I(net_68764),
    .O(net_68805)
  );
  InMux inmux_17_6_68771_68822 (
    .I(net_68771),
    .O(net_68822)
  );
  InMux inmux_17_6_68779_68835 (
    .I(net_68779),
    .O(net_68835)
  );
  InMux inmux_17_6_68783_68827 (
    .I(net_68783),
    .O(net_68827)
  );
  InMux inmux_17_6_68785_68815 (
    .I(net_68785),
    .O(net_68815)
  );
  SRMux inmux_17_6_9_68839 (
    .I(net_9),
    .O(net_68839)
  );
  ClkMux inmux_17_7_5_68961 (
    .I(net_5),
    .O(net_68961)
  );
  InMux inmux_17_7_68888_68958 (
    .I(net_68888),
    .O(net_68958)
  );
  CEMux inmux_17_7_68899_68960 (
    .I(net_68899),
    .O(net_68960)
  );
  SRMux inmux_17_7_9_68962 (
    .I(net_9),
    .O(net_68962)
  );
  ClkMux inmux_17_8_5_69084 (
    .I(net_5),
    .O(net_69084)
  );
  InMux inmux_17_8_69005_69050 (
    .I(net_69005),
    .O(net_69050)
  );
  InMux inmux_17_8_69006_69044 (
    .I(net_69006),
    .O(net_69044)
  );
  InMux inmux_17_8_69009_69043 (
    .I(net_69009),
    .O(net_69043)
  );
  InMux inmux_17_8_69013_69075 (
    .I(net_69013),
    .O(net_69075)
  );
  InMux inmux_17_8_69014_69074 (
    .I(net_69014),
    .O(net_69074)
  );
  InMux inmux_17_8_69019_69051 (
    .I(net_69019),
    .O(net_69051)
  );
  InMux inmux_17_8_69020_69073 (
    .I(net_69020),
    .O(net_69073)
  );
  CEMux inmux_17_8_69022_69083 (
    .I(net_69022),
    .O(net_69083)
  );
  InMux inmux_17_8_69024_69046 (
    .I(net_69024),
    .O(net_69046)
  );
  InMux inmux_17_8_69024_69049 (
    .I(net_69024),
    .O(net_69049)
  );
  InMux inmux_17_8_69028_69045 (
    .I(net_69028),
    .O(net_69045)
  );
  InMux inmux_17_8_69030_69052 (
    .I(net_69030),
    .O(net_69052)
  );
  InMux inmux_17_8_69032_69076 (
    .I(net_69032),
    .O(net_69076)
  );
  ClkMux inmux_17_9_5_69207 (
    .I(net_5),
    .O(net_69207)
  );
  InMux inmux_17_9_69128_69185 (
    .I(net_69128),
    .O(net_69185)
  );
  InMux inmux_17_9_69131_69203 (
    .I(net_69131),
    .O(net_69203)
  );
  SRMux inmux_17_9_9_69208 (
    .I(net_9),
    .O(net_69208)
  );
  IoInMux inmux_18_0_71884_71870 (
    .I(net_71884),
    .O(net_71870)
  );
  ClkMux inmux_18_10_5_73161 (
    .I(net_5),
    .O(net_73161)
  );
  InMux inmux_18_10_73081_73128 (
    .I(net_73081),
    .O(net_73128)
  );
  InMux inmux_18_10_73082_73134 (
    .I(net_73082),
    .O(net_73134)
  );
  InMux inmux_18_10_73086_73146 (
    .I(net_73086),
    .O(net_73146)
  );
  InMux inmux_18_10_73087_73140 (
    .I(net_73087),
    .O(net_73140)
  );
  InMux inmux_18_10_73091_73115 (
    .I(net_73091),
    .O(net_73115)
  );
  InMux inmux_18_10_73094_73116 (
    .I(net_73094),
    .O(net_73116)
  );
  InMux inmux_18_10_73095_73122 (
    .I(net_73095),
    .O(net_73122)
  );
  InMux inmux_18_10_73096_73133 (
    .I(net_73096),
    .O(net_73133)
  );
  InMux inmux_18_10_73097_73121 (
    .I(net_73097),
    .O(net_73121)
  );
  InMux inmux_18_10_73103_73145 (
    .I(net_73103),
    .O(net_73145)
  );
  InMux inmux_18_10_73104_73139 (
    .I(net_73104),
    .O(net_73139)
  );
  InMux inmux_18_10_73106_73157 (
    .I(net_73106),
    .O(net_73157)
  );
  InMux inmux_18_10_73107_73127 (
    .I(net_73107),
    .O(net_73127)
  );
  InMux inmux_18_10_73113_73123 (
    .I(net_73113),
    .O(net_73123)
  );
  InMux inmux_18_10_73119_73129 (
    .I(net_73119),
    .O(net_73129)
  );
  InMux inmux_18_10_73125_73135 (
    .I(net_73125),
    .O(net_73135)
  );
  InMux inmux_18_10_73131_73141 (
    .I(net_73131),
    .O(net_73141)
  );
  InMux inmux_18_10_73137_73147 (
    .I(net_73137),
    .O(net_73147)
  );
  InMux inmux_18_10_73143_73153 (
    .I(net_73143),
    .O(net_73153)
  );
  SRMux inmux_18_10_9_73162 (
    .I(net_9),
    .O(net_73162)
  );
  ClkMux inmux_18_11_5_73284 (
    .I(net_5),
    .O(net_73284)
  );
  InMux inmux_18_11_73205_73250 (
    .I(net_73205),
    .O(net_73250)
  );
  InMux inmux_18_11_73210_73275 (
    .I(net_73210),
    .O(net_73275)
  );
  InMux inmux_18_11_73211_73279 (
    .I(net_73211),
    .O(net_73279)
  );
  InMux inmux_18_11_73218_73243 (
    .I(net_73218),
    .O(net_73243)
  );
  InMux inmux_18_11_73220_73258 (
    .I(net_73220),
    .O(net_73258)
  );
  InMux inmux_18_11_73223_73267 (
    .I(net_73223),
    .O(net_73267)
  );
  InMux inmux_18_11_73225_73240 (
    .I(net_73225),
    .O(net_73240)
  );
  InMux inmux_18_11_73228_73264 (
    .I(net_73228),
    .O(net_73264)
  );
  SRMux inmux_18_11_9_73285 (
    .I(net_9),
    .O(net_73285)
  );
  ClkMux inmux_18_12_5_73407 (
    .I(net_5),
    .O(net_73407)
  );
  InMux inmux_18_12_73330_73375 (
    .I(net_73330),
    .O(net_73375)
  );
  InMux inmux_18_12_73331_73367 (
    .I(net_73331),
    .O(net_73367)
  );
  InMux inmux_18_12_73335_73399 (
    .I(net_73335),
    .O(net_73399)
  );
  InMux inmux_18_12_73336_73381 (
    .I(net_73336),
    .O(net_73381)
  );
  InMux inmux_18_12_73342_73386 (
    .I(net_73342),
    .O(net_73386)
  );
  InMux inmux_18_12_73352_73360 (
    .I(net_73352),
    .O(net_73360)
  );
  InMux inmux_18_12_73353_73404 (
    .I(net_73353),
    .O(net_73404)
  );
  SRMux inmux_18_12_9_73408 (
    .I(net_9),
    .O(net_73408)
  );
  ClkMux inmux_18_13_5_73530 (
    .I(net_5),
    .O(net_73530)
  );
  InMux inmux_18_13_73451_73513 (
    .I(net_73451),
    .O(net_73513)
  );
  InMux inmux_18_13_73459_73507 (
    .I(net_73459),
    .O(net_73507)
  );
  InMux inmux_18_13_73467_73486 (
    .I(net_73467),
    .O(net_73486)
  );
  InMux inmux_18_13_73475_73521 (
    .I(net_73475),
    .O(net_73521)
  );
  InMux inmux_18_13_73477_73497 (
    .I(net_73477),
    .O(net_73497)
  );
  InMux inmux_18_13_73481_73492 (
    .I(net_73481),
    .O(net_73492)
  );
  SRMux inmux_18_13_9_73531 (
    .I(net_9),
    .O(net_73531)
  );
  ClkMux inmux_18_14_5_73653 (
    .I(net_5),
    .O(net_73653)
  );
  InMux inmux_18_14_73573_73608 (
    .I(net_73573),
    .O(net_73608)
  );
  InMux inmux_18_14_73575_73649 (
    .I(net_73575),
    .O(net_73649)
  );
  InMux inmux_18_14_73576_73626 (
    .I(net_73576),
    .O(net_73626)
  );
  InMux inmux_18_14_73582_73618 (
    .I(net_73582),
    .O(net_73618)
  );
  InMux inmux_18_14_73584_73637 (
    .I(net_73584),
    .O(net_73637)
  );
  InMux inmux_18_14_73587_73631 (
    .I(net_73587),
    .O(net_73631)
  );
  InMux inmux_18_14_73590_73612 (
    .I(net_73590),
    .O(net_73612)
  );
  InMux inmux_18_14_73599_73643 (
    .I(net_73599),
    .O(net_73643)
  );
  SRMux inmux_18_14_9_73654 (
    .I(net_9),
    .O(net_73654)
  );
  InMux inmux_18_15_73697_73737 (
    .I(net_73697),
    .O(net_73737)
  );
  InMux inmux_18_15_73698_73767 (
    .I(net_73698),
    .O(net_73767)
  );
  InMux inmux_18_15_73700_73731 (
    .I(net_73700),
    .O(net_73731)
  );
  InMux inmux_18_15_73701_73742 (
    .I(net_73701),
    .O(net_73742)
  );
  InMux inmux_18_15_73702_73760 (
    .I(net_73702),
    .O(net_73760)
  );
  InMux inmux_18_15_73703_73730 (
    .I(net_73703),
    .O(net_73730)
  );
  InMux inmux_18_15_73704_73749 (
    .I(net_73704),
    .O(net_73749)
  );
  InMux inmux_18_15_73705_73743 (
    .I(net_73705),
    .O(net_73743)
  );
  InMux inmux_18_15_73706_73773 (
    .I(net_73706),
    .O(net_73773)
  );
  InMux inmux_18_15_73707_73755 (
    .I(net_73707),
    .O(net_73755)
  );
  InMux inmux_18_15_73708_73761 (
    .I(net_73708),
    .O(net_73761)
  );
  InMux inmux_18_15_73709_73748 (
    .I(net_73709),
    .O(net_73748)
  );
  InMux inmux_18_15_73711_73772 (
    .I(net_73711),
    .O(net_73772)
  );
  InMux inmux_18_15_73722_73766 (
    .I(net_73722),
    .O(net_73766)
  );
  InMux inmux_18_15_73723_73736 (
    .I(net_73723),
    .O(net_73736)
  );
  InMux inmux_18_15_73724_73754 (
    .I(net_73724),
    .O(net_73754)
  );
  InMux inmux_18_15_73728_73738 (
    .I(net_73728),
    .O(net_73738)
  );
  InMux inmux_18_15_73734_73744 (
    .I(net_73734),
    .O(net_73744)
  );
  InMux inmux_18_15_73740_73750 (
    .I(net_73740),
    .O(net_73750)
  );
  InMux inmux_18_15_73746_73756 (
    .I(net_73746),
    .O(net_73756)
  );
  InMux inmux_18_15_73752_73762 (
    .I(net_73752),
    .O(net_73762)
  );
  InMux inmux_18_15_73758_73768 (
    .I(net_73758),
    .O(net_73768)
  );
  InMux inmux_18_15_73764_73774 (
    .I(net_73764),
    .O(net_73774)
  );
  ClkMux inmux_18_16_5_73899 (
    .I(net_5),
    .O(net_73899)
  );
  InMux inmux_18_16_73814_73855 (
    .I(net_73814),
    .O(net_73855)
  );
  InMux inmux_18_16_73819_73859 (
    .I(net_73819),
    .O(net_73859)
  );
  InMux inmux_18_16_73830_73883 (
    .I(net_73830),
    .O(net_73883)
  );
  InMux inmux_18_16_73835_73864 (
    .I(net_73835),
    .O(net_73864)
  );
  InMux inmux_18_16_73839_73876 (
    .I(net_73839),
    .O(net_73876)
  );
  InMux inmux_18_16_73841_73895 (
    .I(net_73841),
    .O(net_73895)
  );
  InMux inmux_18_16_73843_73853 (
    .I(net_73843),
    .O(net_73853)
  );
  InMux inmux_18_16_73844_73852 (
    .I(net_73844),
    .O(net_73852)
  );
  InMux inmux_18_16_73848_73854 (
    .I(net_73848),
    .O(net_73854)
  );
  InMux inmux_18_16_73850_73878 (
    .I(net_73850),
    .O(net_73878)
  );
  SRMux inmux_18_16_9_73900 (
    .I(net_9),
    .O(net_73900)
  );
  ClkMux inmux_18_17_5_74022 (
    .I(net_5),
    .O(net_74022)
  );
  InMux inmux_18_17_73973_73999 (
    .I(net_73973),
    .O(net_73999)
  );
  SRMux inmux_18_17_9_74023 (
    .I(net_9),
    .O(net_74023)
  );
  ClkMux inmux_18_2_5_72177 (
    .I(net_5),
    .O(net_72177)
  );
  InMux inmux_18_2_72103_72154 (
    .I(net_72103),
    .O(net_72154)
  );
  InMux inmux_18_2_72109_72157 (
    .I(net_72109),
    .O(net_72157)
  );
  InMux inmux_18_2_72116_72155 (
    .I(net_72116),
    .O(net_72155)
  );
  SRMux inmux_18_2_9_72178 (
    .I(net_9),
    .O(net_72178)
  );
  IoInMux inmux_18_31_75679_75668 (
    .I(net_75679),
    .O(net_75668)
  );
  IoInMux inmux_18_31_75682_75671 (
    .I(net_75682),
    .O(net_75671)
  );
  ClkMux inmux_18_3_5_72300 (
    .I(net_5),
    .O(net_72300)
  );
  InMux inmux_18_3_72222_72267 (
    .I(net_72222),
    .O(net_72267)
  );
  InMux inmux_18_3_72223_72261 (
    .I(net_72223),
    .O(net_72261)
  );
  InMux inmux_18_3_72224_72272 (
    .I(net_72224),
    .O(net_72272)
  );
  InMux inmux_18_3_72228_72285 (
    .I(net_72228),
    .O(net_72285)
  );
  InMux inmux_18_3_72229_72279 (
    .I(net_72229),
    .O(net_72279)
  );
  InMux inmux_18_3_72233_72253 (
    .I(net_72233),
    .O(net_72253)
  );
  InMux inmux_18_3_72235_72298 (
    .I(net_72235),
    .O(net_72298)
  );
  InMux inmux_18_3_72249_72289 (
    .I(net_72249),
    .O(net_72289)
  );
  SRMux inmux_18_3_9_72301 (
    .I(net_9),
    .O(net_72301)
  );
  InMux inmux_18_4_72344_72420 (
    .I(net_72344),
    .O(net_72420)
  );
  InMux inmux_18_4_72345_72378 (
    .I(net_72345),
    .O(net_72378)
  );
  InMux inmux_18_4_72346_72413 (
    .I(net_72346),
    .O(net_72413)
  );
  InMux inmux_18_4_72347_72395 (
    .I(net_72347),
    .O(net_72395)
  );
  InMux inmux_18_4_72349_72390 (
    .I(net_72349),
    .O(net_72390)
  );
  InMux inmux_18_4_72350_72389 (
    .I(net_72350),
    .O(net_72389)
  );
  InMux inmux_18_4_72351_72384 (
    .I(net_72351),
    .O(net_72384)
  );
  InMux inmux_18_4_72352_72419 (
    .I(net_72352),
    .O(net_72419)
  );
  InMux inmux_18_4_72353_72396 (
    .I(net_72353),
    .O(net_72396)
  );
  InMux inmux_18_4_72354_72407 (
    .I(net_72354),
    .O(net_72407)
  );
  InMux inmux_18_4_72355_72408 (
    .I(net_72355),
    .O(net_72408)
  );
  InMux inmux_18_4_72356_72383 (
    .I(net_72356),
    .O(net_72383)
  );
  InMux inmux_18_4_72358_72402 (
    .I(net_72358),
    .O(net_72402)
  );
  InMux inmux_18_4_72359_72414 (
    .I(net_72359),
    .O(net_72414)
  );
  InMux inmux_18_4_72360_72401 (
    .I(net_72360),
    .O(net_72401)
  );
  InMux inmux_18_4_72364_72377 (
    .I(net_72364),
    .O(net_72377)
  );
  InMux inmux_18_4_72375_72385 (
    .I(net_72375),
    .O(net_72385)
  );
  InMux inmux_18_4_72381_72391 (
    .I(net_72381),
    .O(net_72391)
  );
  InMux inmux_18_4_72387_72397 (
    .I(net_72387),
    .O(net_72397)
  );
  InMux inmux_18_4_72393_72403 (
    .I(net_72393),
    .O(net_72403)
  );
  InMux inmux_18_4_72399_72409 (
    .I(net_72399),
    .O(net_72409)
  );
  InMux inmux_18_4_72405_72415 (
    .I(net_72405),
    .O(net_72415)
  );
  InMux inmux_18_4_72411_72421 (
    .I(net_72411),
    .O(net_72421)
  );
  ClkMux inmux_18_5_5_72546 (
    .I(net_5),
    .O(net_72546)
  );
  InMux inmux_18_5_72461_72502 (
    .I(net_72461),
    .O(net_72502)
  );
  InMux inmux_18_5_72469_72505 (
    .I(net_72469),
    .O(net_72505)
  );
  InMux inmux_18_5_72470_72532 (
    .I(net_72470),
    .O(net_72532)
  );
  InMux inmux_18_5_72472_72506 (
    .I(net_72472),
    .O(net_72506)
  );
  InMux inmux_18_5_72474_72524 (
    .I(net_72474),
    .O(net_72524)
  );
  InMux inmux_18_5_72475_72542 (
    .I(net_72475),
    .O(net_72542)
  );
  InMux inmux_18_5_72477_72511 (
    .I(net_72477),
    .O(net_72511)
  );
  InMux inmux_18_5_72478_72500 (
    .I(net_72478),
    .O(net_72500)
  );
  InMux inmux_18_5_72479_72501 (
    .I(net_72479),
    .O(net_72501)
  );
  InMux inmux_18_5_72482_72537 (
    .I(net_72482),
    .O(net_72537)
  );
  InMux inmux_18_5_72495_72520 (
    .I(net_72495),
    .O(net_72520)
  );
  InMux inmux_18_5_72498_72508 (
    .I(net_72498),
    .O(net_72508)
  );
  SRMux inmux_18_5_9_72547 (
    .I(net_9),
    .O(net_72547)
  );
  ClkMux inmux_18_6_5_72669 (
    .I(net_5),
    .O(net_72669)
  );
  InMux inmux_18_6_72590_72647 (
    .I(net_72590),
    .O(net_72647)
  );
  InMux inmux_18_6_72594_72652 (
    .I(net_72594),
    .O(net_72652)
  );
  InMux inmux_18_6_72597_72642 (
    .I(net_72597),
    .O(net_72642)
  );
  InMux inmux_18_6_72598_72658 (
    .I(net_72598),
    .O(net_72658)
  );
  InMux inmux_18_6_72599_72664 (
    .I(net_72599),
    .O(net_72664)
  );
  InMux inmux_18_6_72604_72624 (
    .I(net_72604),
    .O(net_72624)
  );
  InMux inmux_18_6_72612_72630 (
    .I(net_72612),
    .O(net_72630)
  );
  InMux inmux_18_6_72618_72667 (
    .I(net_72618),
    .O(net_72667)
  );
  SRMux inmux_18_6_9_72670 (
    .I(net_9),
    .O(net_72670)
  );
  ClkMux inmux_18_7_5_72792 (
    .I(net_5),
    .O(net_72792)
  );
  InMux inmux_18_7_72717_72753 (
    .I(net_72717),
    .O(net_72753)
  );
  InMux inmux_18_7_72718_72752 (
    .I(net_72718),
    .O(net_72752)
  );
  InMux inmux_18_7_72719_72746 (
    .I(net_72719),
    .O(net_72746)
  );
  InMux inmux_18_7_72721_72759 (
    .I(net_72721),
    .O(net_72759)
  );
  InMux inmux_18_7_72723_72764 (
    .I(net_72723),
    .O(net_72764)
  );
  InMux inmux_18_7_72725_72771 (
    .I(net_72725),
    .O(net_72771)
  );
  InMux inmux_18_7_72727_72776 (
    .I(net_72727),
    .O(net_72776)
  );
  InMux inmux_18_7_72728_72783 (
    .I(net_72728),
    .O(net_72783)
  );
  InMux inmux_18_7_72730_72788 (
    .I(net_72730),
    .O(net_72788)
  );
  InMux inmux_18_7_72734_72747 (
    .I(net_72734),
    .O(net_72747)
  );
  InMux inmux_18_7_72742_72758 (
    .I(net_72742),
    .O(net_72758)
  );
  InMux inmux_18_7_72742_72765 (
    .I(net_72742),
    .O(net_72765)
  );
  InMux inmux_18_7_72742_72770 (
    .I(net_72742),
    .O(net_72770)
  );
  InMux inmux_18_7_72742_72777 (
    .I(net_72742),
    .O(net_72777)
  );
  InMux inmux_18_7_72742_72782 (
    .I(net_72742),
    .O(net_72782)
  );
  InMux inmux_18_7_72742_72789 (
    .I(net_72742),
    .O(net_72789)
  );
  InMux inmux_18_7_72744_72754 (
    .I(net_72744),
    .O(net_72754)
  );
  InMux inmux_18_7_72750_72760 (
    .I(net_72750),
    .O(net_72760)
  );
  InMux inmux_18_7_72756_72766 (
    .I(net_72756),
    .O(net_72766)
  );
  InMux inmux_18_7_72762_72772 (
    .I(net_72762),
    .O(net_72772)
  );
  InMux inmux_18_7_72768_72778 (
    .I(net_72768),
    .O(net_72778)
  );
  InMux inmux_18_7_72774_72784 (
    .I(net_72774),
    .O(net_72784)
  );
  InMux inmux_18_7_72780_72790 (
    .I(net_72780),
    .O(net_72790)
  );
  SRMux inmux_18_7_9_72793 (
    .I(net_9),
    .O(net_72793)
  );
  ClkMux inmux_18_8_5_72915 (
    .I(net_5),
    .O(net_72915)
  );
  InMux inmux_18_8_72830_72871 (
    .I(net_72830),
    .O(net_72871)
  );
  InMux inmux_18_8_72836_72893 (
    .I(net_72836),
    .O(net_72893)
  );
  InMux inmux_18_8_72840_72898 (
    .I(net_72840),
    .O(net_72898)
  );
  InMux inmux_18_8_72846_72870 (
    .I(net_72846),
    .O(net_72870)
  );
  InMux inmux_18_8_72848_72913 (
    .I(net_72848),
    .O(net_72913)
  );
  InMux inmux_18_8_72850_72875 (
    .I(net_72850),
    .O(net_72875)
  );
  InMux inmux_18_8_72854_72869 (
    .I(net_72854),
    .O(net_72869)
  );
  InMux inmux_18_8_72854_72874 (
    .I(net_72854),
    .O(net_72874)
  );
  InMux inmux_18_8_72867_72877 (
    .I(net_72867),
    .O(net_72877)
  );
  SRMux inmux_18_8_9_72916 (
    .I(net_9),
    .O(net_72916)
  );
  ClkMux inmux_18_9_5_73038 (
    .I(net_5),
    .O(net_73038)
  );
  InMux inmux_18_9_72970_72997 (
    .I(net_72970),
    .O(net_72997)
  );
  InMux inmux_18_9_72971_73022 (
    .I(net_72971),
    .O(net_73022)
  );
  InMux inmux_18_9_72973_73029 (
    .I(net_72973),
    .O(net_73029)
  );
  InMux inmux_18_9_72974_73012 (
    .I(net_72974),
    .O(net_73012)
  );
  InMux inmux_18_9_72976_72993 (
    .I(net_72976),
    .O(net_72993)
  );
  InMux inmux_18_9_72987_72991 (
    .I(net_72987),
    .O(net_72991)
  );
  SRMux inmux_18_9_9_73039 (
    .I(net_9),
    .O(net_73039)
  );
  ClkMux inmux_1_10_5_8158 (
    .I(net_5),
    .O(net_8158)
  );
  InMux inmux_1_10_8081_8143 (
    .I(net_8081),
    .O(net_8143)
  );
  InMux inmux_1_10_8083_8124 (
    .I(net_8083),
    .O(net_8124)
  );
  InMux inmux_1_10_8085_8136 (
    .I(net_8085),
    .O(net_8136)
  );
  InMux inmux_1_10_8089_8120 (
    .I(net_8089),
    .O(net_8120)
  );
  InMux inmux_1_10_8095_8131 (
    .I(net_8095),
    .O(net_8131)
  );
  InMux inmux_1_10_8098_8149 (
    .I(net_8098),
    .O(net_8149)
  );
  InMux inmux_1_10_8104_8114 (
    .I(net_8104),
    .O(net_8114)
  );
  InMux inmux_1_10_8108_8155 (
    .I(net_8108),
    .O(net_8155)
  );
  SRMux inmux_1_10_9_8159 (
    .I(net_9),
    .O(net_8159)
  );
  ClkMux inmux_1_11_5_8305 (
    .I(net_5),
    .O(net_8305)
  );
  InMux inmux_1_11_8228_8283 (
    .I(net_8228),
    .O(net_8283)
  );
  InMux inmux_1_11_8232_8271 (
    .I(net_8232),
    .O(net_8271)
  );
  InMux inmux_1_11_8235_8276 (
    .I(net_8235),
    .O(net_8276)
  );
  InMux inmux_1_11_8246_8266 (
    .I(net_8246),
    .O(net_8266)
  );
  InMux inmux_1_11_8247_8294 (
    .I(net_8247),
    .O(net_8294)
  );
  InMux inmux_1_11_8248_8261 (
    .I(net_8248),
    .O(net_8261)
  );
  InMux inmux_1_11_8252_8303 (
    .I(net_8252),
    .O(net_8303)
  );
  InMux inmux_1_11_8254_8291 (
    .I(net_8254),
    .O(net_8291)
  );
  SRMux inmux_1_11_9_8306 (
    .I(net_9),
    .O(net_8306)
  );
  ClkMux inmux_1_12_5_8452 (
    .I(net_5),
    .O(net_8452)
  );
  InMux inmux_1_12_8375_8430 (
    .I(net_8375),
    .O(net_8430)
  );
  InMux inmux_1_12_8377_8418 (
    .I(net_8377),
    .O(net_8418)
  );
  InMux inmux_1_12_8378_8424 (
    .I(net_8378),
    .O(net_8424)
  );
  InMux inmux_1_12_8380_8444 (
    .I(net_8380),
    .O(net_8444)
  );
  InMux inmux_1_12_8383_8450 (
    .I(net_8383),
    .O(net_8450)
  );
  InMux inmux_1_12_8384_8406 (
    .I(net_8384),
    .O(net_8406)
  );
  InMux inmux_1_12_8392_8438 (
    .I(net_8392),
    .O(net_8438)
  );
  SRMux inmux_1_12_9_8453 (
    .I(net_9),
    .O(net_8453)
  );
  ClkMux inmux_1_13_5_8599 (
    .I(net_5),
    .O(net_8599)
  );
  InMux inmux_1_13_8519_8564 (
    .I(net_8519),
    .O(net_8564)
  );
  InMux inmux_1_13_8522_8582 (
    .I(net_8522),
    .O(net_8582)
  );
  InMux inmux_1_13_8525_8573 (
    .I(net_8525),
    .O(net_8573)
  );
  InMux inmux_1_13_8527_8560 (
    .I(net_8527),
    .O(net_8560)
  );
  InMux inmux_1_13_8529_8591 (
    .I(net_8529),
    .O(net_8591)
  );
  InMux inmux_1_13_8531_8594 (
    .I(net_8531),
    .O(net_8594)
  );
  InMux inmux_1_13_8533_8553 (
    .I(net_8533),
    .O(net_8553)
  );
  InMux inmux_1_13_8535_8576 (
    .I(net_8535),
    .O(net_8576)
  );
  SRMux inmux_1_13_9_8600 (
    .I(net_9),
    .O(net_8600)
  );
  ClkMux inmux_1_14_5_8746 (
    .I(net_5),
    .O(net_8746)
  );
  InMux inmux_1_14_8669_8719 (
    .I(net_8669),
    .O(net_8719)
  );
  InMux inmux_1_14_8670_8735 (
    .I(net_8670),
    .O(net_8735)
  );
  InMux inmux_1_14_8671_8726 (
    .I(net_8671),
    .O(net_8726)
  );
  InMux inmux_1_14_8673_8707 (
    .I(net_8673),
    .O(net_8707)
  );
  InMux inmux_1_14_8680_8714 (
    .I(net_8680),
    .O(net_8714)
  );
  InMux inmux_1_14_8683_8743 (
    .I(net_8683),
    .O(net_8743)
  );
  InMux inmux_1_14_8684_8730 (
    .I(net_8684),
    .O(net_8730)
  );
  InMux inmux_1_14_8689_8700 (
    .I(net_8689),
    .O(net_8700)
  );
  SRMux inmux_1_14_9_8747 (
    .I(net_9),
    .O(net_8747)
  );
  ClkMux inmux_1_15_5_8893 (
    .I(net_5),
    .O(net_8893)
  );
  InMux inmux_1_15_8813_8882 (
    .I(net_8813),
    .O(net_8882)
  );
  InMux inmux_1_15_8824_8879 (
    .I(net_8824),
    .O(net_8879)
  );
  InMux inmux_1_15_8827_8861 (
    .I(net_8827),
    .O(net_8861)
  );
  InMux inmux_1_15_8829_8891 (
    .I(net_8829),
    .O(net_8891)
  );
  InMux inmux_1_15_8830_8866 (
    .I(net_8830),
    .O(net_8866)
  );
  InMux inmux_1_15_8835_8870 (
    .I(net_8835),
    .O(net_8870)
  );
  InMux inmux_1_15_8838_8846 (
    .I(net_8838),
    .O(net_8846)
  );
  InMux inmux_1_15_8841_8854 (
    .I(net_8841),
    .O(net_8854)
  );
  SRMux inmux_1_15_9_8894 (
    .I(net_9),
    .O(net_8894)
  );
  ClkMux inmux_1_16_5_9040 (
    .I(net_5),
    .O(net_9040)
  );
  InMux inmux_1_16_8965_8996 (
    .I(net_8965),
    .O(net_8996)
  );
  InMux inmux_1_16_8977_9001 (
    .I(net_8977),
    .O(net_9001)
  );
  InMux inmux_1_16_8981_9008 (
    .I(net_8981),
    .O(net_9008)
  );
  InMux inmux_1_16_8982_9014 (
    .I(net_8982),
    .O(net_9014)
  );
  InMux inmux_1_16_8984_9018 (
    .I(net_8984),
    .O(net_9018)
  );
  InMux inmux_1_16_8988_9030 (
    .I(net_8988),
    .O(net_9030)
  );
  InMux inmux_1_16_8989_9024 (
    .I(net_8989),
    .O(net_9024)
  );
  SRMux inmux_1_16_9_9041 (
    .I(net_9),
    .O(net_9041)
  );
  ClkMux inmux_1_17_5_9187 (
    .I(net_5),
    .O(net_9187)
  );
  InMux inmux_1_17_9107_9159 (
    .I(net_9107),
    .O(net_9159)
  );
  InMux inmux_1_17_9108_9146 (
    .I(net_9108),
    .O(net_9146)
  );
  InMux inmux_1_17_9111_9154 (
    .I(net_9111),
    .O(net_9154)
  );
  InMux inmux_1_17_9130_9182 (
    .I(net_9130),
    .O(net_9182)
  );
  SRMux inmux_1_17_9_9188 (
    .I(net_9),
    .O(net_9188)
  );
  ClkMux inmux_1_18_5_9334 (
    .I(net_5),
    .O(net_9334)
  );
  InMux inmux_1_18_9256_9289 (
    .I(net_9256),
    .O(net_9289)
  );
  InMux inmux_1_18_9261_9295 (
    .I(net_9261),
    .O(net_9295)
  );
  InMux inmux_1_18_9267_9311 (
    .I(net_9267),
    .O(net_9311)
  );
  InMux inmux_1_18_9281_9323 (
    .I(net_9281),
    .O(net_9323)
  );
  SRMux inmux_1_18_9_9335 (
    .I(net_9),
    .O(net_9335)
  );
  ClkMux inmux_1_19_5_9481 (
    .I(net_5),
    .O(net_9481)
  );
  InMux inmux_1_19_9402_9476 (
    .I(net_9402),
    .O(net_9476)
  );
  InMux inmux_1_19_9407_9436 (
    .I(net_9407),
    .O(net_9436)
  );
  InMux inmux_1_19_9416_9465 (
    .I(net_9416),
    .O(net_9465)
  );
  SRMux inmux_1_19_9_9482 (
    .I(net_9),
    .O(net_9482)
  );
  ClkMux inmux_1_1_5_6795 (
    .I(net_5),
    .O(net_6795)
  );
  InMux inmux_1_1_6717_6784 (
    .I(net_6717),
    .O(net_6784)
  );
  InMux inmux_1_1_6720_6792 (
    .I(net_6720),
    .O(net_6792)
  );
  InMux inmux_1_1_6721_6779 (
    .I(net_6721),
    .O(net_6779)
  );
  InMux inmux_1_1_6726_6760 (
    .I(net_6726),
    .O(net_6760)
  );
  InMux inmux_1_1_6727_6763 (
    .I(net_6727),
    .O(net_6763)
  );
  InMux inmux_1_1_6727_6778 (
    .I(net_6727),
    .O(net_6778)
  );
  InMux inmux_1_1_6730_6781 (
    .I(net_6730),
    .O(net_6781)
  );
  InMux inmux_1_1_6745_6761 (
    .I(net_6745),
    .O(net_6761)
  );
  SRMux inmux_1_1_9_6796 (
    .I(net_9),
    .O(net_6796)
  );
  ClkMux inmux_1_20_5_9628 (
    .I(net_5),
    .O(net_9628)
  );
  InMux inmux_1_20_9554_9617 (
    .I(net_9554),
    .O(net_9617)
  );
  InMux inmux_1_20_9560_9596 (
    .I(net_9560),
    .O(net_9596)
  );
  InMux inmux_1_20_9564_9590 (
    .I(net_9564),
    .O(net_9590)
  );
  InMux inmux_1_20_9576_9625 (
    .I(net_9576),
    .O(net_9625)
  );
  SRMux inmux_1_20_9_9629 (
    .I(net_9),
    .O(net_9629)
  );
  ClkMux inmux_1_21_5_9775 (
    .I(net_5),
    .O(net_9775)
  );
  InMux inmux_1_21_9700_9748 (
    .I(net_9700),
    .O(net_9748)
  );
  InMux inmux_1_21_9721_9729 (
    .I(net_9721),
    .O(net_9729)
  );
  SRMux inmux_1_21_9_9776 (
    .I(net_9),
    .O(net_9776)
  );
  ClkMux inmux_1_22_5_9922 (
    .I(net_5),
    .O(net_9922)
  );
  InMux inmux_1_22_9843_9905 (
    .I(net_9843),
    .O(net_9905)
  );
  InMux inmux_1_22_9848_9913 (
    .I(net_9848),
    .O(net_9913)
  );
  InMux inmux_1_22_9851_9882 (
    .I(net_9851),
    .O(net_9882)
  );
  SRMux inmux_1_22_9_9923 (
    .I(net_9),
    .O(net_9923)
  );
  InMux inmux_1_23_10015_10037 (
    .I(net_10015),
    .O(net_10037)
  );
  ClkMux inmux_1_23_5_10069 (
    .I(net_5),
    .O(net_10069)
  );
  SRMux inmux_1_23_9_10070 (
    .I(net_9),
    .O(net_10070)
  );
  ClkMux inmux_1_2_5_6982 (
    .I(net_5),
    .O(net_6982)
  );
  InMux inmux_1_2_6904_6978 (
    .I(net_6904),
    .O(net_6978)
  );
  InMux inmux_1_2_6905_6977 (
    .I(net_6905),
    .O(net_6977)
  );
  InMux inmux_1_2_6907_6979 (
    .I(net_6907),
    .O(net_6979)
  );
  InMux inmux_1_2_6909_6967 (
    .I(net_6909),
    .O(net_6967)
  );
  InMux inmux_1_2_6912_6955 (
    .I(net_6912),
    .O(net_6955)
  );
  InMux inmux_1_2_6915_6971 (
    .I(net_6915),
    .O(net_6971)
  );
  InMux inmux_1_2_6917_6937 (
    .I(net_6917),
    .O(net_6937)
  );
  InMux inmux_1_2_6917_6944 (
    .I(net_6917),
    .O(net_6944)
  );
  InMux inmux_1_2_6919_6960 (
    .I(net_6919),
    .O(net_6960)
  );
  InMux inmux_1_2_6922_6980 (
    .I(net_6922),
    .O(net_6980)
  );
  InMux inmux_1_2_6924_6949 (
    .I(net_6924),
    .O(net_6949)
  );
  InMux inmux_1_2_6925_6943 (
    .I(net_6925),
    .O(net_6943)
  );
  InMux inmux_1_2_6940_6950 (
    .I(net_6940),
    .O(net_6950)
  );
  InMux inmux_1_2_6946_6956 (
    .I(net_6946),
    .O(net_6956)
  );
  InMux inmux_1_2_6952_6962 (
    .I(net_6952),
    .O(net_6962)
  );
  InMux inmux_1_2_6958_6968 (
    .I(net_6958),
    .O(net_6968)
  );
  InMux inmux_1_2_6964_6974 (
    .I(net_6964),
    .O(net_6974)
  );
  SRMux inmux_1_2_9_6983 (
    .I(net_9),
    .O(net_6983)
  );
  ClkMux inmux_1_3_5_7129 (
    .I(net_5),
    .O(net_7129)
  );
  InMux inmux_1_3_7050_7090 (
    .I(net_7050),
    .O(net_7090)
  );
  InMux inmux_1_3_7050_7119 (
    .I(net_7050),
    .O(net_7119)
  );
  InMux inmux_1_3_7052_7124 (
    .I(net_7052),
    .O(net_7124)
  );
  InMux inmux_1_3_7056_7126 (
    .I(net_7056),
    .O(net_7126)
  );
  InMux inmux_1_3_7057_7121 (
    .I(net_7057),
    .O(net_7121)
  );
  InMux inmux_1_3_7058_7108 (
    .I(net_7058),
    .O(net_7108)
  );
  InMux inmux_1_3_7060_7082 (
    .I(net_7060),
    .O(net_7082)
  );
  InMux inmux_1_3_7060_7118 (
    .I(net_7060),
    .O(net_7118)
  );
  InMux inmux_1_3_7062_7127 (
    .I(net_7062),
    .O(net_7127)
  );
  InMux inmux_1_3_7065_7096 (
    .I(net_7065),
    .O(net_7096)
  );
  InMux inmux_1_3_7066_7114 (
    .I(net_7066),
    .O(net_7114)
  );
  InMux inmux_1_3_7072_7100 (
    .I(net_7072),
    .O(net_7100)
  );
  InMux inmux_1_3_7074_7084 (
    .I(net_7074),
    .O(net_7084)
  );
  InMux inmux_1_3_7074_7089 (
    .I(net_7074),
    .O(net_7089)
  );
  InMux inmux_1_3_7075_7085 (
    .I(net_7075),
    .O(net_7085)
  );
  InMux inmux_1_3_7077_7088 (
    .I(net_7077),
    .O(net_7088)
  );
  InMux inmux_1_3_7078_7120 (
    .I(net_7078),
    .O(net_7120)
  );
  SRMux inmux_1_3_9_7130 (
    .I(net_9),
    .O(net_7130)
  );
  ClkMux inmux_1_4_5_7276 (
    .I(net_5),
    .O(net_7276)
  );
  InMux inmux_1_4_7196_7248 (
    .I(net_7196),
    .O(net_7248)
  );
  InMux inmux_1_4_7199_7271 (
    .I(net_7199),
    .O(net_7271)
  );
  InMux inmux_1_4_7201_7273 (
    .I(net_7201),
    .O(net_7273)
  );
  InMux inmux_1_4_7205_7236 (
    .I(net_7205),
    .O(net_7236)
  );
  InMux inmux_1_4_7207_7272 (
    .I(net_7207),
    .O(net_7272)
  );
  InMux inmux_1_4_7209_7265 (
    .I(net_7209),
    .O(net_7265)
  );
  InMux inmux_1_4_7213_7254 (
    .I(net_7213),
    .O(net_7254)
  );
  InMux inmux_1_4_7214_7231 (
    .I(net_7214),
    .O(net_7231)
  );
  InMux inmux_1_4_7214_7238 (
    .I(net_7214),
    .O(net_7238)
  );
  InMux inmux_1_4_7218_7274 (
    .I(net_7218),
    .O(net_7274)
  );
  InMux inmux_1_4_7222_7242 (
    .I(net_7222),
    .O(net_7242)
  );
  InMux inmux_1_4_7226_7261 (
    .I(net_7226),
    .O(net_7261)
  );
  InMux inmux_1_4_7234_7244 (
    .I(net_7234),
    .O(net_7244)
  );
  InMux inmux_1_4_7240_7250 (
    .I(net_7240),
    .O(net_7250)
  );
  InMux inmux_1_4_7246_7256 (
    .I(net_7246),
    .O(net_7256)
  );
  InMux inmux_1_4_7252_7262 (
    .I(net_7252),
    .O(net_7262)
  );
  InMux inmux_1_4_7258_7268 (
    .I(net_7258),
    .O(net_7268)
  );
  SRMux inmux_1_4_9_7277 (
    .I(net_9),
    .O(net_7277)
  );
  ClkMux inmux_1_5_5_7423 (
    .I(net_5),
    .O(net_7423)
  );
  InMux inmux_1_5_7343_7407 (
    .I(net_7343),
    .O(net_7407)
  );
  InMux inmux_1_5_7346_7415 (
    .I(net_7346),
    .O(net_7415)
  );
  InMux inmux_1_5_7349_7402 (
    .I(net_7349),
    .O(net_7402)
  );
  InMux inmux_1_5_7353_7418 (
    .I(net_7353),
    .O(net_7418)
  );
  InMux inmux_1_5_7357_7408 (
    .I(net_7357),
    .O(net_7408)
  );
  InMux inmux_1_5_7359_7409 (
    .I(net_7359),
    .O(net_7409)
  );
  InMux inmux_1_5_7361_7390 (
    .I(net_7361),
    .O(net_7390)
  );
  InMux inmux_1_5_7363_7395 (
    .I(net_7363),
    .O(net_7395)
  );
  InMux inmux_1_5_7364_7377 (
    .I(net_7364),
    .O(net_7377)
  );
  InMux inmux_1_5_7366_7384 (
    .I(net_7366),
    .O(net_7384)
  );
  SRMux inmux_1_5_9_7424 (
    .I(net_9),
    .O(net_7424)
  );
  ClkMux inmux_1_6_5_7570 (
    .I(net_5),
    .O(net_7570)
  );
  InMux inmux_1_6_7491_7543 (
    .I(net_7491),
    .O(net_7543)
  );
  InMux inmux_1_6_7506_7549 (
    .I(net_7506),
    .O(net_7549)
  );
  InMux inmux_1_6_7509_7529 (
    .I(net_7509),
    .O(net_7529)
  );
  InMux inmux_1_6_7510_7554 (
    .I(net_7510),
    .O(net_7554)
  );
  InMux inmux_1_6_7519_7561 (
    .I(net_7519),
    .O(net_7561)
  );
  SRMux inmux_1_6_9_7571 (
    .I(net_9),
    .O(net_7571)
  );
  ClkMux inmux_1_7_5_7717 (
    .I(net_5),
    .O(net_7717)
  );
  CEMux inmux_1_7_7648_7716 (
    .I(net_7648),
    .O(net_7716)
  );
  InMux inmux_1_7_7651_7676 (
    .I(net_7651),
    .O(net_7676)
  );
  ClkMux inmux_1_8_5_7864 (
    .I(net_5),
    .O(net_7864)
  );
  InMux inmux_1_8_7792_7842 (
    .I(net_7792),
    .O(net_7842)
  );
  InMux inmux_1_8_7798_7861 (
    .I(net_7798),
    .O(net_7861)
  );
  InMux inmux_1_8_7801_7835 (
    .I(net_7801),
    .O(net_7835)
  );
  InMux inmux_1_8_7802_7853 (
    .I(net_7802),
    .O(net_7853)
  );
  InMux inmux_1_8_7806_7850 (
    .I(net_7806),
    .O(net_7850)
  );
  InMux inmux_1_8_7808_7823 (
    .I(net_7808),
    .O(net_7823)
  );
  InMux inmux_1_8_7812_7832 (
    .I(net_7812),
    .O(net_7832)
  );
  InMux inmux_1_8_7815_7817 (
    .I(net_7815),
    .O(net_7817)
  );
  SRMux inmux_1_8_9_7865 (
    .I(net_9),
    .O(net_7865)
  );
  ClkMux inmux_1_9_5_8011 (
    .I(net_5),
    .O(net_8011)
  );
  InMux inmux_1_9_7931_8007 (
    .I(net_7931),
    .O(net_8007)
  );
  InMux inmux_1_9_7936_7982 (
    .I(net_7936),
    .O(net_7982)
  );
  InMux inmux_1_9_7944_7973 (
    .I(net_7944),
    .O(net_7973)
  );
  InMux inmux_1_9_7946_7966 (
    .I(net_7946),
    .O(net_7966)
  );
  InMux inmux_1_9_7956_8000 (
    .I(net_7956),
    .O(net_8000)
  );
  InMux inmux_1_9_7960_7997 (
    .I(net_7960),
    .O(net_7997)
  );
  InMux inmux_1_9_7961_7977 (
    .I(net_7961),
    .O(net_7977)
  );
  InMux inmux_1_9_7962_7988 (
    .I(net_7962),
    .O(net_7988)
  );
  SRMux inmux_1_9_9_8012 (
    .I(net_9),
    .O(net_8012)
  );
  ClkMux inmux_20_10_5_80192 (
    .I(net_5),
    .O(net_80192)
  );
  InMux inmux_20_10_80113_80146 (
    .I(net_80113),
    .O(net_80146)
  );
  InMux inmux_20_10_80113_80151 (
    .I(net_80113),
    .O(net_80151)
  );
  InMux inmux_20_10_80113_80170 (
    .I(net_80113),
    .O(net_80170)
  );
  InMux inmux_20_10_80113_80175 (
    .I(net_80113),
    .O(net_80175)
  );
  CEMux inmux_20_10_80114_80191 (
    .I(net_80114),
    .O(net_80191)
  );
  InMux inmux_20_10_80118_80152 (
    .I(net_80118),
    .O(net_80152)
  );
  InMux inmux_20_10_80119_80177 (
    .I(net_80119),
    .O(net_80177)
  );
  InMux inmux_20_10_80126_80148 (
    .I(net_80126),
    .O(net_80148)
  );
  InMux inmux_20_10_80127_80169 (
    .I(net_80127),
    .O(net_80169)
  );
  SRMux inmux_20_10_9_80193 (
    .I(net_9),
    .O(net_80193)
  );
  ClkMux inmux_20_11_5_80315 (
    .I(net_5),
    .O(net_80315)
  );
  InMux inmux_20_11_80242_80307 (
    .I(net_80242),
    .O(net_80307)
  );
  InMux inmux_20_11_80244_80311 (
    .I(net_80244),
    .O(net_80311)
  );
  SRMux inmux_20_11_9_80316 (
    .I(net_9),
    .O(net_80316)
  );
  ClkMux inmux_20_12_5_80438 (
    .I(net_5),
    .O(net_80438)
  );
  CEMux inmux_20_12_6_80437 (
    .I(net_6),
    .O(net_80437)
  );
  InMux inmux_20_12_80362_80405 (
    .I(net_80362),
    .O(net_80405)
  );
  InMux inmux_20_12_80383_80403 (
    .I(net_80383),
    .O(net_80403)
  );
  SRMux inmux_20_12_9_80439 (
    .I(net_9),
    .O(net_80439)
  );
  ClkMux inmux_20_14_5_80684 (
    .I(net_5),
    .O(net_80684)
  );
  CEMux inmux_20_14_80615_80683 (
    .I(net_80615),
    .O(net_80683)
  );
  InMux inmux_20_14_80631_80658 (
    .I(net_80631),
    .O(net_80658)
  );
  ClkMux inmux_20_2_5_79208 (
    .I(net_5),
    .O(net_79208)
  );
  InMux inmux_20_2_79130_79173 (
    .I(net_79130),
    .O(net_79173)
  );
  InMux inmux_20_2_79130_79204 (
    .I(net_79130),
    .O(net_79204)
  );
  InMux inmux_20_2_79143_79175 (
    .I(net_79143),
    .O(net_79175)
  );
  InMux inmux_20_2_79143_79206 (
    .I(net_79143),
    .O(net_79206)
  );
  CEMux inmux_20_2_79155_79207 (
    .I(net_79155),
    .O(net_79207)
  );
  SRMux inmux_20_2_9_79209 (
    .I(net_9),
    .O(net_79209)
  );
  ClkMux inmux_20_3_5_79331 (
    .I(net_5),
    .O(net_79331)
  );
  InMux inmux_20_3_79259_79326 (
    .I(net_79259),
    .O(net_79326)
  );
  InMux inmux_20_3_79260_79293 (
    .I(net_79260),
    .O(net_79293)
  );
  InMux inmux_20_3_79268_79314 (
    .I(net_79268),
    .O(net_79314)
  );
  InMux inmux_20_3_79270_79302 (
    .I(net_79270),
    .O(net_79302)
  );
  InMux inmux_20_3_79278_79320 (
    .I(net_79278),
    .O(net_79320)
  );
  InMux inmux_20_3_79279_79287 (
    .I(net_79279),
    .O(net_79287)
  );
  SRMux inmux_20_3_9_79332 (
    .I(net_9),
    .O(net_79332)
  );
  ClkMux inmux_20_4_5_79454 (
    .I(net_5),
    .O(net_79454)
  );
  InMux inmux_20_4_79387_79414 (
    .I(net_79387),
    .O(net_79414)
  );
  InMux inmux_20_4_79388_79415 (
    .I(net_79388),
    .O(net_79415)
  );
  CEMux inmux_20_4_79401_79453 (
    .I(net_79401),
    .O(net_79453)
  );
  SRMux inmux_20_4_9_79455 (
    .I(net_9),
    .O(net_79455)
  );
  ClkMux inmux_20_5_5_79577 (
    .I(net_5),
    .O(net_79577)
  );
  InMux inmux_20_5_79501_79530 (
    .I(net_79501),
    .O(net_79530)
  );
  InMux inmux_20_5_79504_79543 (
    .I(net_79504),
    .O(net_79543)
  );
  InMux inmux_20_5_79505_79538 (
    .I(net_79505),
    .O(net_79538)
  );
  InMux inmux_20_5_79508_79563 (
    .I(net_79508),
    .O(net_79563)
  );
  InMux inmux_20_5_79519_79573 (
    .I(net_79519),
    .O(net_79573)
  );
  InMux inmux_20_5_79522_79551 (
    .I(net_79522),
    .O(net_79551)
  );
  InMux inmux_20_5_79527_79569 (
    .I(net_79527),
    .O(net_79569)
  );
  InMux inmux_20_5_79528_79554 (
    .I(net_79528),
    .O(net_79554)
  );
  SRMux inmux_20_5_9_79578 (
    .I(net_9),
    .O(net_79578)
  );
  ClkMux inmux_20_6_5_79700 (
    .I(net_5),
    .O(net_79700)
  );
  InMux inmux_20_6_79630_79678 (
    .I(net_79630),
    .O(net_79678)
  );
  InMux inmux_20_6_79631_79684 (
    .I(net_79631),
    .O(net_79684)
  );
  InMux inmux_20_6_79632_79654 (
    .I(net_79632),
    .O(net_79654)
  );
  InMux inmux_20_6_79632_79680 (
    .I(net_79632),
    .O(net_79680)
  );
  InMux inmux_20_6_79632_79685 (
    .I(net_79632),
    .O(net_79685)
  );
  InMux inmux_20_6_79633_79653 (
    .I(net_79633),
    .O(net_79653)
  );
  InMux inmux_20_6_79640_79677 (
    .I(net_79640),
    .O(net_79677)
  );
  InMux inmux_20_6_79641_79683 (
    .I(net_79641),
    .O(net_79683)
  );
  InMux inmux_20_6_79642_79686 (
    .I(net_79642),
    .O(net_79686)
  );
  InMux inmux_20_6_79645_79679 (
    .I(net_79645),
    .O(net_79679)
  );
  InMux inmux_20_6_79646_79656 (
    .I(net_79646),
    .O(net_79656)
  );
  CEMux inmux_20_6_79647_79699 (
    .I(net_79647),
    .O(net_79699)
  );
  InMux inmux_20_6_79649_79655 (
    .I(net_79649),
    .O(net_79655)
  );
  SRMux inmux_20_6_9_79701 (
    .I(net_9),
    .O(net_79701)
  );
  ClkMux inmux_20_7_5_79823 (
    .I(net_5),
    .O(net_79823)
  );
  CEMux inmux_20_7_79745_79822 (
    .I(net_79745),
    .O(net_79822)
  );
  InMux inmux_20_7_79750_79808 (
    .I(net_79750),
    .O(net_79808)
  );
  InMux inmux_20_7_79752_79809 (
    .I(net_79752),
    .O(net_79809)
  );
  InMux inmux_20_7_79757_79806 (
    .I(net_79757),
    .O(net_79806)
  );
  InMux inmux_20_7_79770_79807 (
    .I(net_79770),
    .O(net_79807)
  );
  SRMux inmux_20_7_9_79824 (
    .I(net_9),
    .O(net_79824)
  );
  ClkMux inmux_20_8_5_79946 (
    .I(net_5),
    .O(net_79946)
  );
  InMux inmux_20_8_79893_79937 (
    .I(net_79893),
    .O(net_79937)
  );
  SRMux inmux_20_8_9_79947 (
    .I(net_9),
    .O(net_79947)
  );
  ClkMux inmux_20_9_5_80069 (
    .I(net_5),
    .O(net_80069)
  );
  InMux inmux_20_9_79996_80066 (
    .I(net_79996),
    .O(net_80066)
  );
  InMux inmux_20_9_79998_80043 (
    .I(net_79998),
    .O(net_80043)
  );
  InMux inmux_20_9_80004_80048 (
    .I(net_80004),
    .O(net_80048)
  );
  InMux inmux_20_9_80020_80053 (
    .I(net_80020),
    .O(net_80053)
  );
  SRMux inmux_20_9_9_80070 (
    .I(net_9),
    .O(net_80070)
  );
  IoInMux inmux_21_0_82750_82732 (
    .I(net_82750),
    .O(net_82732)
  );
  ClkMux inmux_21_10_5_84023 (
    .I(net_5),
    .O(net_84023)
  );
  InMux inmux_21_10_83943_83983 (
    .I(net_83943),
    .O(net_83983)
  );
  InMux inmux_21_10_83951_84001 (
    .I(net_83951),
    .O(net_84001)
  );
  InMux inmux_21_10_83954_83995 (
    .I(net_83954),
    .O(net_83995)
  );
  InMux inmux_21_10_83956_83976 (
    .I(net_83956),
    .O(net_83976)
  );
  InMux inmux_21_10_83958_83990 (
    .I(net_83958),
    .O(net_83990)
  );
  SRMux inmux_21_10_9_84024 (
    .I(net_9),
    .O(net_84024)
  );
  ClkMux inmux_21_3_5_83162 (
    .I(net_5),
    .O(net_83162)
  );
  InMux inmux_21_3_83100_83115 (
    .I(net_83100),
    .O(net_83115)
  );
  InMux inmux_21_3_83102_83134 (
    .I(net_83102),
    .O(net_83134)
  );
  InMux inmux_21_3_83106_83130 (
    .I(net_83106),
    .O(net_83130)
  );
  InMux inmux_21_3_83112_83157 (
    .I(net_83112),
    .O(net_83157)
  );
  SRMux inmux_21_3_9_83163 (
    .I(net_9),
    .O(net_83163)
  );
  ClkMux inmux_21_4_5_83285 (
    .I(net_5),
    .O(net_83285)
  );
  InMux inmux_21_4_83206_83270 (
    .I(net_83206),
    .O(net_83270)
  );
  InMux inmux_21_4_83219_83244 (
    .I(net_83219),
    .O(net_83244)
  );
  InMux inmux_21_4_83227_83252 (
    .I(net_83227),
    .O(net_83252)
  );
  InMux inmux_21_4_83228_83280 (
    .I(net_83228),
    .O(net_83280)
  );
  InMux inmux_21_4_83236_83238 (
    .I(net_83236),
    .O(net_83238)
  );
  SRMux inmux_21_4_9_83286 (
    .I(net_9),
    .O(net_83286)
  );
  ClkMux inmux_21_5_5_83408 (
    .I(net_5),
    .O(net_83408)
  );
  InMux inmux_21_5_83328_83385 (
    .I(net_83328),
    .O(net_83385)
  );
  InMux inmux_21_5_83356_83376 (
    .I(net_83356),
    .O(net_83376)
  );
  InMux inmux_21_5_83357_83399 (
    .I(net_83357),
    .O(net_83399)
  );
  SRMux inmux_21_5_9_83409 (
    .I(net_9),
    .O(net_83409)
  );
  ClkMux inmux_21_6_5_83531 (
    .I(net_5),
    .O(net_83531)
  );
  InMux inmux_21_6_83452_83526 (
    .I(net_83452),
    .O(net_83526)
  );
  InMux inmux_21_6_83471_83522 (
    .I(net_83471),
    .O(net_83522)
  );
  InMux inmux_21_6_83479_83514 (
    .I(net_83479),
    .O(net_83514)
  );
  InMux inmux_21_6_83481_83509 (
    .I(net_83481),
    .O(net_83509)
  );
  SRMux inmux_21_6_9_83532 (
    .I(net_9),
    .O(net_83532)
  );
  ClkMux inmux_21_7_5_83654 (
    .I(net_5),
    .O(net_83654)
  );
  InMux inmux_21_7_83576_83614 (
    .I(net_83576),
    .O(net_83614)
  );
  InMux inmux_21_7_83577_83622 (
    .I(net_83577),
    .O(net_83622)
  );
  InMux inmux_21_7_83579_83649 (
    .I(net_83579),
    .O(net_83649)
  );
  InMux inmux_21_7_83600_83627 (
    .I(net_83600),
    .O(net_83627)
  );
  SRMux inmux_21_7_9_83655 (
    .I(net_9),
    .O(net_83655)
  );
  ClkMux inmux_21_8_5_83777 (
    .I(net_5),
    .O(net_83777)
  );
  InMux inmux_21_8_83699_83737 (
    .I(net_83699),
    .O(net_83737)
  );
  InMux inmux_21_8_83701_83744 (
    .I(net_83701),
    .O(net_83744)
  );
  InMux inmux_21_8_83703_83756 (
    .I(net_83703),
    .O(net_83756)
  );
  InMux inmux_21_8_83704_83774 (
    .I(net_83704),
    .O(net_83774)
  );
  InMux inmux_21_8_83706_83749 (
    .I(net_83706),
    .O(net_83749)
  );
  InMux inmux_21_8_83707_83755 (
    .I(net_83707),
    .O(net_83755)
  );
  InMux inmux_21_8_83710_83761 (
    .I(net_83710),
    .O(net_83761)
  );
  InMux inmux_21_8_83711_83731 (
    .I(net_83711),
    .O(net_83731)
  );
  InMux inmux_21_8_83716_83743 (
    .I(net_83716),
    .O(net_83743)
  );
  InMux inmux_21_8_83717_83768 (
    .I(net_83717),
    .O(net_83768)
  );
  InMux inmux_21_8_83719_83773 (
    .I(net_83719),
    .O(net_83773)
  );
  InMux inmux_21_8_83720_83767 (
    .I(net_83720),
    .O(net_83767)
  );
  InMux inmux_21_8_83721_83738 (
    .I(net_83721),
    .O(net_83738)
  );
  InMux inmux_21_8_83725_83750 (
    .I(net_83725),
    .O(net_83750)
  );
  InMux inmux_21_8_83726_83732 (
    .I(net_83726),
    .O(net_83732)
  );
  InMux inmux_21_8_83727_83762 (
    .I(net_83727),
    .O(net_83762)
  );
  InMux inmux_21_8_83729_83739 (
    .I(net_83729),
    .O(net_83739)
  );
  InMux inmux_21_8_83735_83745 (
    .I(net_83735),
    .O(net_83745)
  );
  InMux inmux_21_8_83741_83751 (
    .I(net_83741),
    .O(net_83751)
  );
  InMux inmux_21_8_83747_83757 (
    .I(net_83747),
    .O(net_83757)
  );
  InMux inmux_21_8_83753_83763 (
    .I(net_83753),
    .O(net_83763)
  );
  InMux inmux_21_8_83759_83769 (
    .I(net_83759),
    .O(net_83769)
  );
  InMux inmux_21_8_83765_83775 (
    .I(net_83765),
    .O(net_83775)
  );
  SRMux inmux_21_8_9_83778 (
    .I(net_9),
    .O(net_83778)
  );
  ClkMux inmux_21_9_5_83900 (
    .I(net_5),
    .O(net_83900)
  );
  InMux inmux_21_9_83815_83856 (
    .I(net_83815),
    .O(net_83856)
  );
  InMux inmux_21_9_83825_83897 (
    .I(net_83825),
    .O(net_83897)
  );
  InMux inmux_21_9_83830_83861 (
    .I(net_83830),
    .O(net_83861)
  );
  InMux inmux_21_9_83831_83855 (
    .I(net_83831),
    .O(net_83855)
  );
  InMux inmux_21_9_83832_83866 (
    .I(net_83832),
    .O(net_83866)
  );
  InMux inmux_21_9_83834_83854 (
    .I(net_83834),
    .O(net_83854)
  );
  InMux inmux_21_9_83835_83889 (
    .I(net_83835),
    .O(net_83889)
  );
  InMux inmux_21_9_83836_83860 (
    .I(net_83836),
    .O(net_83860)
  );
  InMux inmux_21_9_83840_83877 (
    .I(net_83840),
    .O(net_83877)
  );
  InMux inmux_21_9_83847_83867 (
    .I(net_83847),
    .O(net_83867)
  );
  InMux inmux_21_9_83850_83895 (
    .I(net_83850),
    .O(net_83895)
  );
  InMux inmux_21_9_83852_83862 (
    .I(net_83852),
    .O(net_83862)
  );
  InMux inmux_21_9_83858_83868 (
    .I(net_83858),
    .O(net_83868)
  );
  InMux inmux_21_9_83864_83874 (
    .I(net_83864),
    .O(net_83874)
  );
  SRMux inmux_21_9_9_83901 (
    .I(net_9),
    .O(net_83901)
  );
  IoInMux inmux_22_0_86583_86563 (
    .I(net_86583),
    .O(net_86563)
  );
  ClkMux inmux_22_3_5_86993 (
    .I(net_5),
    .O(net_86993)
  );
  InMux inmux_22_3_86917_86972 (
    .I(net_86917),
    .O(net_86972)
  );
  InMux inmux_22_3_86924_86960 (
    .I(net_86924),
    .O(net_86960)
  );
  InMux inmux_22_3_86940_86948 (
    .I(net_86940),
    .O(net_86948)
  );
  SRMux inmux_22_3_9_86994 (
    .I(net_9),
    .O(net_86994)
  );
  ClkMux inmux_22_4_5_87116 (
    .I(net_5),
    .O(net_87116)
  );
  InMux inmux_22_4_87036_87105 (
    .I(net_87036),
    .O(net_87105)
  );
  InMux inmux_22_4_87054_87083 (
    .I(net_87054),
    .O(net_87083)
  );
  InMux inmux_22_4_87059_87113 (
    .I(net_87059),
    .O(net_87113)
  );
  SRMux inmux_22_4_9_87117 (
    .I(net_9),
    .O(net_87117)
  );
  ClkMux inmux_22_5_5_87239 (
    .I(net_5),
    .O(net_87239)
  );
  InMux inmux_22_5_87163_87218 (
    .I(net_87163),
    .O(net_87218)
  );
  InMux inmux_22_5_87176_87210 (
    .I(net_87176),
    .O(net_87210)
  );
  InMux inmux_22_5_87177_87192 (
    .I(net_87177),
    .O(net_87192)
  );
  InMux inmux_22_5_87178_87236 (
    .I(net_87178),
    .O(net_87236)
  );
  InMux inmux_22_5_87183_87231 (
    .I(net_87183),
    .O(net_87231)
  );
  SRMux inmux_22_5_9_87240 (
    .I(net_9),
    .O(net_87240)
  );
  ClkMux inmux_22_6_5_87362 (
    .I(net_5),
    .O(net_87362)
  );
  InMux inmux_22_6_87301_87342 (
    .I(net_87301),
    .O(net_87342)
  );
  InMux inmux_22_6_87305_87354 (
    .I(net_87305),
    .O(net_87354)
  );
  SRMux inmux_22_6_9_87363 (
    .I(net_9),
    .O(net_87363)
  );
  ClkMux inmux_22_7_5_87485 (
    .I(net_5),
    .O(net_87485)
  );
  InMux inmux_22_7_87413_87453 (
    .I(net_87413),
    .O(net_87453)
  );
  InMux inmux_22_7_87428_87465 (
    .I(net_87428),
    .O(net_87465)
  );
  InMux inmux_22_7_87430_87469 (
    .I(net_87430),
    .O(net_87469)
  );
  InMux inmux_22_7_87434_87483 (
    .I(net_87434),
    .O(net_87483)
  );
  SRMux inmux_22_7_9_87486 (
    .I(net_9),
    .O(net_87486)
  );
  ClkMux inmux_22_8_5_87608 (
    .I(net_5),
    .O(net_87608)
  );
  InMux inmux_22_8_87539_87563 (
    .I(net_87539),
    .O(net_87563)
  );
  InMux inmux_22_8_87542_87588 (
    .I(net_87542),
    .O(net_87588)
  );
  InMux inmux_22_8_87543_87575 (
    .I(net_87543),
    .O(net_87575)
  );
  InMux inmux_22_8_87547_87600 (
    .I(net_87547),
    .O(net_87600)
  );
  InMux inmux_22_8_87550_87582 (
    .I(net_87550),
    .O(net_87582)
  );
  InMux inmux_22_8_87557_87594 (
    .I(net_87557),
    .O(net_87594)
  );
  SRMux inmux_22_8_9_87609 (
    .I(net_9),
    .O(net_87609)
  );
  ClkMux inmux_22_9_5_87731 (
    .I(net_5),
    .O(net_87731)
  );
  InMux inmux_22_9_87665_87709 (
    .I(net_87665),
    .O(net_87709)
  );
  InMux inmux_22_9_87668_87702 (
    .I(net_87668),
    .O(net_87702)
  );
  InMux inmux_22_9_87676_87727 (
    .I(net_87676),
    .O(net_87727)
  );
  InMux inmux_22_9_87677_87721 (
    .I(net_87677),
    .O(net_87721)
  );
  InMux inmux_22_9_87682_87684 (
    .I(net_87682),
    .O(net_87684)
  );
  SRMux inmux_22_9_9_87732 (
    .I(net_9),
    .O(net_87732)
  );
  IoInMux inmux_23_0_90410_90394 (
    .I(net_90410),
    .O(net_90394)
  );
  ClkMux inmux_23_5_5_91070 (
    .I(net_5),
    .O(net_91070)
  );
  InMux inmux_23_5_90991_91053 (
    .I(net_90991),
    .O(net_91053)
  );
  InMux inmux_23_5_91009_91067 (
    .I(net_91009),
    .O(net_91067)
  );
  InMux inmux_23_5_91014_91048 (
    .I(net_91014),
    .O(net_91048)
  );
  InMux inmux_23_5_91018_91031 (
    .I(net_91018),
    .O(net_91031)
  );
  InMux inmux_23_5_91021_91023 (
    .I(net_91021),
    .O(net_91023)
  );
  SRMux inmux_23_5_9_91071 (
    .I(net_9),
    .O(net_91071)
  );
  ClkMux inmux_23_6_5_91193 (
    .I(net_5),
    .O(net_91193)
  );
  InMux inmux_23_6_91133_91165 (
    .I(net_91133),
    .O(net_91165)
  );
  InMux inmux_23_6_91137_91152 (
    .I(net_91137),
    .O(net_91152)
  );
  InMux inmux_23_6_91141_91188 (
    .I(net_91141),
    .O(net_91188)
  );
  SRMux inmux_23_6_9_91194 (
    .I(net_9),
    .O(net_91194)
  );
  ClkMux inmux_23_8_5_91439 (
    .I(net_5),
    .O(net_91439)
  );
  InMux inmux_23_8_91380_91434 (
    .I(net_91380),
    .O(net_91434)
  );
  SRMux inmux_23_8_9_91440 (
    .I(net_9),
    .O(net_91440)
  );
  ClkMux inmux_23_9_5_91562 (
    .I(net_5),
    .O(net_91562)
  );
  InMux inmux_23_9_91495_91536 (
    .I(net_91495),
    .O(net_91536)
  );
  SRMux inmux_23_9_9_91563 (
    .I(net_9),
    .O(net_91563)
  );
  InMux inmux_25_11_100150_100197 (
    .I(net_100150),
    .O(net_100197)
  );
  InMux inmux_25_11_100154_100194 (
    .I(net_100154),
    .O(net_100194)
  );
  InMux inmux_25_11_100155_100195 (
    .I(net_100155),
    .O(net_100195)
  );
  InMux inmux_25_11_100156_100185 (
    .I(net_100156),
    .O(net_100185)
  );
  InMux inmux_25_11_100164_100183 (
    .I(net_100164),
    .O(net_100183)
  );
  InMux inmux_25_11_100168_100186 (
    .I(net_100168),
    .O(net_100186)
  );
  InMux inmux_25_11_100169_100184 (
    .I(net_100169),
    .O(net_100184)
  );
  InMux inmux_25_11_100170_100190 (
    .I(net_100170),
    .O(net_100190)
  );
  InMux inmux_25_11_100171_100187 (
    .I(net_100171),
    .O(net_100187)
  );
  InMux inmux_25_11_100172_100193 (
    .I(net_100172),
    .O(net_100193)
  );
  InMux inmux_25_11_100173_100188 (
    .I(net_100173),
    .O(net_100188)
  );
  InMux inmux_25_11_100175_100189 (
    .I(net_100175),
    .O(net_100189)
  );
  InMux inmux_25_11_100176_100196 (
    .I(net_100176),
    .O(net_100196)
  );
  InMux inmux_25_11_100178_100191 (
    .I(net_100178),
    .O(net_100191)
  );
  InMux inmux_25_11_100180_100192 (
    .I(net_100180),
    .O(net_100192)
  );
  InMux inmux_25_11_100181_100198 (
    .I(net_100181),
    .O(net_100198)
  );
  InMux inmux_25_12_100302_100347 (
    .I(net_100302),
    .O(net_100347)
  );
  InMux inmux_25_12_100303_100333 (
    .I(net_100303),
    .O(net_100333)
  );
  InMux inmux_25_12_100309_100340 (
    .I(net_100309),
    .O(net_100340)
  );
  InMux inmux_25_12_100310_100338 (
    .I(net_100310),
    .O(net_100338)
  );
  InMux inmux_25_12_100311_100343 (
    .I(net_100311),
    .O(net_100343)
  );
  InMux inmux_25_12_100312_100345 (
    .I(net_100312),
    .O(net_100345)
  );
  InMux inmux_25_12_100313_100335 (
    .I(net_100313),
    .O(net_100335)
  );
  InMux inmux_25_12_100314_100334 (
    .I(net_100314),
    .O(net_100334)
  );
  InMux inmux_25_12_100317_100341 (
    .I(net_100317),
    .O(net_100341)
  );
  InMux inmux_25_12_100318_100348 (
    .I(net_100318),
    .O(net_100348)
  );
  InMux inmux_25_12_100319_100342 (
    .I(net_100319),
    .O(net_100342)
  );
  InMux inmux_25_12_100320_100344 (
    .I(net_100320),
    .O(net_100344)
  );
  InMux inmux_25_12_100325_100336 (
    .I(net_100325),
    .O(net_100336)
  );
  InMux inmux_25_12_100326_100346 (
    .I(net_100326),
    .O(net_100346)
  );
  InMux inmux_25_12_100330_100337 (
    .I(net_100330),
    .O(net_100337)
  );
  InMux inmux_25_12_100331_100339 (
    .I(net_100331),
    .O(net_100339)
  );
  InMux inmux_25_6_99370_99409 (
    .I(net_99370),
    .O(net_99409)
  );
  InMux inmux_25_6_99373_99412 (
    .I(net_99373),
    .O(net_99412)
  );
  InMux inmux_25_6_99380_99411 (
    .I(net_99380),
    .O(net_99411)
  );
  InMux inmux_25_6_99383_99405 (
    .I(net_99383),
    .O(net_99405)
  );
  InMux inmux_25_6_99385_99413 (
    .I(net_99385),
    .O(net_99413)
  );
  InMux inmux_25_6_99386_99417 (
    .I(net_99386),
    .O(net_99417)
  );
  InMux inmux_25_6_99388_99418 (
    .I(net_99388),
    .O(net_99418)
  );
  InMux inmux_25_6_99389_99403 (
    .I(net_99389),
    .O(net_99403)
  );
  InMux inmux_25_6_99391_99408 (
    .I(net_99391),
    .O(net_99408)
  );
  InMux inmux_25_6_99394_99407 (
    .I(net_99394),
    .O(net_99407)
  );
  InMux inmux_25_6_99395_99414 (
    .I(net_99395),
    .O(net_99414)
  );
  InMux inmux_25_6_99396_99415 (
    .I(net_99396),
    .O(net_99415)
  );
  InMux inmux_25_6_99398_99416 (
    .I(net_99398),
    .O(net_99416)
  );
  InMux inmux_25_6_99399_99406 (
    .I(net_99399),
    .O(net_99406)
  );
  InMux inmux_25_6_99400_99404 (
    .I(net_99400),
    .O(net_99404)
  );
  InMux inmux_25_6_99401_99410 (
    .I(net_99401),
    .O(net_99410)
  );
  InMux inmux_25_7_99520_99567 (
    .I(net_99520),
    .O(net_99567)
  );
  InMux inmux_25_7_99521_99553 (
    .I(net_99521),
    .O(net_99553)
  );
  InMux inmux_25_7_99523_99566 (
    .I(net_99523),
    .O(net_99566)
  );
  InMux inmux_25_7_99527_99557 (
    .I(net_99527),
    .O(net_99557)
  );
  InMux inmux_25_7_99529_99563 (
    .I(net_99529),
    .O(net_99563)
  );
  InMux inmux_25_7_99530_99565 (
    .I(net_99530),
    .O(net_99565)
  );
  InMux inmux_25_7_99532_99561 (
    .I(net_99532),
    .O(net_99561)
  );
  InMux inmux_25_7_99533_99555 (
    .I(net_99533),
    .O(net_99555)
  );
  InMux inmux_25_7_99534_99562 (
    .I(net_99534),
    .O(net_99562)
  );
  InMux inmux_25_7_99535_99568 (
    .I(net_99535),
    .O(net_99568)
  );
  InMux inmux_25_7_99536_99556 (
    .I(net_99536),
    .O(net_99556)
  );
  InMux inmux_25_7_99543_99554 (
    .I(net_99543),
    .O(net_99554)
  );
  InMux inmux_25_7_99544_99558 (
    .I(net_99544),
    .O(net_99558)
  );
  InMux inmux_25_7_99545_99559 (
    .I(net_99545),
    .O(net_99559)
  );
  InMux inmux_25_7_99547_99564 (
    .I(net_99547),
    .O(net_99564)
  );
  InMux inmux_25_7_99549_99560 (
    .I(net_99549),
    .O(net_99560)
  );
  CEMux inmux_2_10_10_12497 (
    .I(net_10),
    .O(net_12497)
  );
  InMux inmux_2_10_12419_12476 (
    .I(net_12419),
    .O(net_12476)
  );
  InMux inmux_2_10_12432_12483 (
    .I(net_12432),
    .O(net_12483)
  );
  InMux inmux_2_10_12433_12477 (
    .I(net_12433),
    .O(net_12477)
  );
  InMux inmux_2_10_12436_12475 (
    .I(net_12436),
    .O(net_12475)
  );
  InMux inmux_2_10_12439_12488 (
    .I(net_12439),
    .O(net_12488)
  );
  InMux inmux_2_10_12442_12452 (
    .I(net_12442),
    .O(net_12452)
  );
  InMux inmux_2_10_12443_12496 (
    .I(net_12443),
    .O(net_12496)
  );
  InMux inmux_2_10_12446_12464 (
    .I(net_12446),
    .O(net_12464)
  );
  ClkMux inmux_2_10_5_12498 (
    .I(net_5),
    .O(net_12498)
  );
  InMux inmux_2_11_12541_12617 (
    .I(net_12541),
    .O(net_12617)
  );
  InMux inmux_2_11_12542_12587 (
    .I(net_12542),
    .O(net_12587)
  );
  InMux inmux_2_11_12544_12594 (
    .I(net_12544),
    .O(net_12594)
  );
  InMux inmux_2_11_12546_12611 (
    .I(net_12546),
    .O(net_12611)
  );
  InMux inmux_2_11_12553_12575 (
    .I(net_12553),
    .O(net_12575)
  );
  InMux inmux_2_11_12554_12600 (
    .I(net_12554),
    .O(net_12600)
  );
  InMux inmux_2_11_12556_12576 (
    .I(net_12556),
    .O(net_12576)
  );
  InMux inmux_2_11_12559_12588 (
    .I(net_12559),
    .O(net_12588)
  );
  InMux inmux_2_11_12563_12612 (
    .I(net_12563),
    .O(net_12612)
  );
  InMux inmux_2_11_12564_12618 (
    .I(net_12564),
    .O(net_12618)
  );
  InMux inmux_2_11_12565_12606 (
    .I(net_12565),
    .O(net_12606)
  );
  InMux inmux_2_11_12566_12581 (
    .I(net_12566),
    .O(net_12581)
  );
  InMux inmux_2_11_12567_12582 (
    .I(net_12567),
    .O(net_12582)
  );
  InMux inmux_2_11_12568_12593 (
    .I(net_12568),
    .O(net_12593)
  );
  InMux inmux_2_11_12569_12599 (
    .I(net_12569),
    .O(net_12599)
  );
  InMux inmux_2_11_12570_12605 (
    .I(net_12570),
    .O(net_12605)
  );
  InMux inmux_2_11_12573_12583 (
    .I(net_12573),
    .O(net_12583)
  );
  InMux inmux_2_11_12579_12589 (
    .I(net_12579),
    .O(net_12589)
  );
  InMux inmux_2_11_12585_12595 (
    .I(net_12585),
    .O(net_12595)
  );
  InMux inmux_2_11_12591_12601 (
    .I(net_12591),
    .O(net_12601)
  );
  InMux inmux_2_11_12597_12607 (
    .I(net_12597),
    .O(net_12607)
  );
  InMux inmux_2_11_12603_12613 (
    .I(net_12603),
    .O(net_12613)
  );
  InMux inmux_2_11_12609_12619 (
    .I(net_12609),
    .O(net_12619)
  );
  ClkMux inmux_2_11_5_12621 (
    .I(net_5),
    .O(net_12621)
  );
  SRMux inmux_2_11_9_12622 (
    .I(net_9),
    .O(net_12622)
  );
  InMux inmux_2_12_12659_12700 (
    .I(net_12659),
    .O(net_12700)
  );
  InMux inmux_2_12_12667_12717 (
    .I(net_12667),
    .O(net_12717)
  );
  InMux inmux_2_12_12669_12722 (
    .I(net_12669),
    .O(net_12722)
  );
  InMux inmux_2_12_12681_12741 (
    .I(net_12681),
    .O(net_12741)
  );
  InMux inmux_2_12_12683_12710 (
    .I(net_12683),
    .O(net_12710)
  );
  InMux inmux_2_12_12685_12729 (
    .I(net_12685),
    .O(net_12729)
  );
  InMux inmux_2_12_12688_12705 (
    .I(net_12688),
    .O(net_12705)
  );
  InMux inmux_2_12_12690_12734 (
    .I(net_12690),
    .O(net_12734)
  );
  InMux inmux_2_12_12692_12698 (
    .I(net_12692),
    .O(net_12698)
  );
  InMux inmux_2_12_12695_12699 (
    .I(net_12695),
    .O(net_12699)
  );
  InMux inmux_2_12_12695_12704 (
    .I(net_12695),
    .O(net_12704)
  );
  InMux inmux_2_12_12695_12711 (
    .I(net_12695),
    .O(net_12711)
  );
  InMux inmux_2_12_12695_12716 (
    .I(net_12695),
    .O(net_12716)
  );
  InMux inmux_2_12_12695_12723 (
    .I(net_12695),
    .O(net_12723)
  );
  InMux inmux_2_12_12695_12728 (
    .I(net_12695),
    .O(net_12728)
  );
  InMux inmux_2_12_12695_12735 (
    .I(net_12695),
    .O(net_12735)
  );
  InMux inmux_2_12_12695_12740 (
    .I(net_12695),
    .O(net_12740)
  );
  InMux inmux_2_12_12696_12706 (
    .I(net_12696),
    .O(net_12706)
  );
  InMux inmux_2_12_12702_12712 (
    .I(net_12702),
    .O(net_12712)
  );
  InMux inmux_2_12_12708_12718 (
    .I(net_12708),
    .O(net_12718)
  );
  InMux inmux_2_12_12714_12724 (
    .I(net_12714),
    .O(net_12724)
  );
  InMux inmux_2_12_12720_12730 (
    .I(net_12720),
    .O(net_12730)
  );
  InMux inmux_2_12_12726_12736 (
    .I(net_12726),
    .O(net_12736)
  );
  InMux inmux_2_12_12732_12742 (
    .I(net_12732),
    .O(net_12742)
  );
  ClkMux inmux_2_12_5_12744 (
    .I(net_5),
    .O(net_12744)
  );
  SRMux inmux_2_12_9_12745 (
    .I(net_9),
    .O(net_12745)
  );
  InMux inmux_2_13_12782_12823 (
    .I(net_12782),
    .O(net_12823)
  );
  InMux inmux_2_13_12790_12840 (
    .I(net_12790),
    .O(net_12840)
  );
  InMux inmux_2_13_12793_12820 (
    .I(net_12793),
    .O(net_12820)
  );
  InMux inmux_2_13_12798_12832 (
    .I(net_12798),
    .O(net_12832)
  );
  InMux inmux_2_13_12802_12822 (
    .I(net_12802),
    .O(net_12822)
  );
  InMux inmux_2_13_12804_12857 (
    .I(net_12804),
    .O(net_12857)
  );
  InMux inmux_2_13_12810_12828 (
    .I(net_12810),
    .O(net_12828)
  );
  InMux inmux_2_13_12812_12853 (
    .I(net_12812),
    .O(net_12853)
  );
  InMux inmux_2_13_12814_12844 (
    .I(net_12814),
    .O(net_12844)
  );
  InMux inmux_2_13_12816_12865 (
    .I(net_12816),
    .O(net_12865)
  );
  InMux inmux_2_13_12818_12863 (
    .I(net_12818),
    .O(net_12863)
  );
  ClkMux inmux_2_13_5_12867 (
    .I(net_5),
    .O(net_12867)
  );
  SRMux inmux_2_13_9_12868 (
    .I(net_9),
    .O(net_12868)
  );
  InMux inmux_2_14_12913_12944 (
    .I(net_12913),
    .O(net_12944)
  );
  InMux inmux_2_14_12913_12982 (
    .I(net_12913),
    .O(net_12982)
  );
  InMux inmux_2_14_12919_12950 (
    .I(net_12919),
    .O(net_12950)
  );
  InMux inmux_2_14_12920_12956 (
    .I(net_12920),
    .O(net_12956)
  );
  InMux inmux_2_14_12925_12945 (
    .I(net_12925),
    .O(net_12945)
  );
  InMux inmux_2_14_12925_12979 (
    .I(net_12925),
    .O(net_12979)
  );
  InMux inmux_2_14_12927_12985 (
    .I(net_12927),
    .O(net_12985)
  );
  InMux inmux_2_14_12928_12962 (
    .I(net_12928),
    .O(net_12962)
  );
  InMux inmux_2_14_12931_12975 (
    .I(net_12931),
    .O(net_12975)
  );
  InMux inmux_2_14_12932_12967 (
    .I(net_12932),
    .O(net_12967)
  );
  InMux inmux_2_14_12934_12951 (
    .I(net_12934),
    .O(net_12951)
  );
  InMux inmux_2_14_12935_12957 (
    .I(net_12935),
    .O(net_12957)
  );
  InMux inmux_2_14_12942_12952 (
    .I(net_12942),
    .O(net_12952)
  );
  InMux inmux_2_14_12948_12958 (
    .I(net_12948),
    .O(net_12958)
  );
  ClkMux inmux_2_14_5_12990 (
    .I(net_5),
    .O(net_12990)
  );
  SRMux inmux_2_14_9_12991 (
    .I(net_9),
    .O(net_12991)
  );
  InMux inmux_2_15_13034_13079 (
    .I(net_13034),
    .O(net_13079)
  );
  InMux inmux_2_15_13035_13068 (
    .I(net_13035),
    .O(net_13068)
  );
  InMux inmux_2_15_13035_13085 (
    .I(net_13035),
    .O(net_13085)
  );
  InMux inmux_2_15_13036_13086 (
    .I(net_13036),
    .O(net_13086)
  );
  InMux inmux_2_15_13037_13111 (
    .I(net_13037),
    .O(net_13111)
  );
  InMux inmux_2_15_13039_13073 (
    .I(net_13039),
    .O(net_13073)
  );
  InMux inmux_2_15_13040_13067 (
    .I(net_13040),
    .O(net_13067)
  );
  InMux inmux_2_15_13040_13084 (
    .I(net_13040),
    .O(net_13084)
  );
  InMux inmux_2_15_13043_13074 (
    .I(net_13043),
    .O(net_13074)
  );
  InMux inmux_2_15_13055_13097 (
    .I(net_13055),
    .O(net_13097)
  );
  InMux inmux_2_15_13060_13080 (
    .I(net_13060),
    .O(net_13080)
  );
  InMux inmux_2_15_13062_13090 (
    .I(net_13062),
    .O(net_13090)
  );
  InMux inmux_2_15_13063_13105 (
    .I(net_13063),
    .O(net_13105)
  );
  InMux inmux_2_15_13065_13075 (
    .I(net_13065),
    .O(net_13075)
  );
  InMux inmux_2_15_13071_13081 (
    .I(net_13071),
    .O(net_13081)
  );
  ClkMux inmux_2_15_5_13113 (
    .I(net_5),
    .O(net_13113)
  );
  SRMux inmux_2_15_9_13114 (
    .I(net_9),
    .O(net_13114)
  );
  InMux inmux_2_16_13158_13189 (
    .I(net_13158),
    .O(net_13189)
  );
  InMux inmux_2_16_13163_13214 (
    .I(net_13163),
    .O(net_13214)
  );
  InMux inmux_2_16_13164_13207 (
    .I(net_13164),
    .O(net_13207)
  );
  InMux inmux_2_16_13166_13233 (
    .I(net_13166),
    .O(net_13233)
  );
  InMux inmux_2_16_13173_13219 (
    .I(net_13173),
    .O(net_13219)
  );
  InMux inmux_2_16_13174_13227 (
    .I(net_13174),
    .O(net_13227)
  );
  InMux inmux_2_16_13183_13198 (
    .I(net_13183),
    .O(net_13198)
  );
  InMux inmux_2_16_13187_13203 (
    .I(net_13187),
    .O(net_13203)
  );
  ClkMux inmux_2_16_5_13236 (
    .I(net_5),
    .O(net_13236)
  );
  SRMux inmux_2_16_9_13237 (
    .I(net_9),
    .O(net_13237)
  );
  InMux inmux_2_17_13291_13356 (
    .I(net_13291),
    .O(net_13356)
  );
  InMux inmux_2_17_13294_13345 (
    .I(net_13294),
    .O(net_13345)
  );
  InMux inmux_2_17_13301_13324 (
    .I(net_13301),
    .O(net_13324)
  );
  ClkMux inmux_2_17_5_13359 (
    .I(net_5),
    .O(net_13359)
  );
  SRMux inmux_2_17_9_13360 (
    .I(net_9),
    .O(net_13360)
  );
  InMux inmux_2_18_13403_13472 (
    .I(net_13403),
    .O(net_13472)
  );
  InMux inmux_2_18_13407_13479 (
    .I(net_13407),
    .O(net_13479)
  );
  InMux inmux_2_18_13408_13444 (
    .I(net_13408),
    .O(net_13444)
  );
  InMux inmux_2_18_13409_13460 (
    .I(net_13409),
    .O(net_13460)
  );
  InMux inmux_2_18_13421_13436 (
    .I(net_13421),
    .O(net_13436)
  );
  ClkMux inmux_2_18_5_13482 (
    .I(net_5),
    .O(net_13482)
  );
  SRMux inmux_2_18_9_13483 (
    .I(net_9),
    .O(net_13483)
  );
  InMux inmux_2_19_13528_13576 (
    .I(net_13528),
    .O(net_13576)
  );
  InMux inmux_2_19_13529_13596 (
    .I(net_13529),
    .O(net_13596)
  );
  InMux inmux_2_19_13531_13560 (
    .I(net_13531),
    .O(net_13560)
  );
  InMux inmux_2_19_13533_13583 (
    .I(net_13533),
    .O(net_13583)
  );
  InMux inmux_2_19_13537_13600 (
    .I(net_13537),
    .O(net_13600)
  );
  InMux inmux_2_19_13538_13567 (
    .I(net_13538),
    .O(net_13567)
  );
  InMux inmux_2_19_13540_13591 (
    .I(net_13540),
    .O(net_13591)
  );
  ClkMux inmux_2_19_5_13605 (
    .I(net_5),
    .O(net_13605)
  );
  SRMux inmux_2_19_9_13606 (
    .I(net_9),
    .O(net_13606)
  );
  InMux inmux_2_1_11272_11305 (
    .I(net_11272),
    .O(net_11305)
  );
  InMux inmux_2_1_11272_11346 (
    .I(net_11272),
    .O(net_11346)
  );
  InMux inmux_2_1_11278_11322 (
    .I(net_11278),
    .O(net_11322)
  );
  InMux inmux_2_1_11279_11324 (
    .I(net_11279),
    .O(net_11324)
  );
  InMux inmux_2_1_11283_11307 (
    .I(net_11283),
    .O(net_11307)
  );
  InMux inmux_2_1_11293_11304 (
    .I(net_11293),
    .O(net_11304)
  );
  InMux inmux_2_1_11293_11325 (
    .I(net_11293),
    .O(net_11325)
  );
  InMux inmux_2_1_11294_11348 (
    .I(net_11294),
    .O(net_11348)
  );
  InMux inmux_2_1_11295_11310 (
    .I(net_11295),
    .O(net_11310)
  );
  InMux inmux_2_1_11295_11336 (
    .I(net_11295),
    .O(net_11336)
  );
  InMux inmux_2_1_11302_11323 (
    .I(net_11302),
    .O(net_11323)
  );
  ClkMux inmux_2_1_5_11351 (
    .I(net_5),
    .O(net_11351)
  );
  SRMux inmux_2_1_9_11352 (
    .I(net_9),
    .O(net_11352)
  );
  InMux inmux_2_20_13650_13690 (
    .I(net_13650),
    .O(net_13690)
  );
  InMux inmux_2_20_13652_13700 (
    .I(net_13652),
    .O(net_13700)
  );
  InMux inmux_2_20_13653_13708 (
    .I(net_13653),
    .O(net_13708)
  );
  InMux inmux_2_20_13655_13711 (
    .I(net_13655),
    .O(net_13711)
  );
  InMux inmux_2_20_13672_13723 (
    .I(net_13672),
    .O(net_13723)
  );
  ClkMux inmux_2_20_5_13728 (
    .I(net_5),
    .O(net_13728)
  );
  SRMux inmux_2_20_9_13729 (
    .I(net_9),
    .O(net_13729)
  );
  InMux inmux_2_21_13776_13829 (
    .I(net_13776),
    .O(net_13829)
  );
  InMux inmux_2_21_13779_13810 (
    .I(net_13779),
    .O(net_13810)
  );
  ClkMux inmux_2_21_5_13851 (
    .I(net_5),
    .O(net_13851)
  );
  SRMux inmux_2_21_9_13852 (
    .I(net_9),
    .O(net_13852)
  );
  InMux inmux_2_22_13897_13959 (
    .I(net_13897),
    .O(net_13959)
  );
  InMux inmux_2_22_13920_13928 (
    .I(net_13920),
    .O(net_13928)
  );
  ClkMux inmux_2_22_5_13974 (
    .I(net_5),
    .O(net_13974)
  );
  SRMux inmux_2_22_9_13975 (
    .I(net_9),
    .O(net_13975)
  );
  InMux inmux_2_23_14026_14074 (
    .I(net_14026),
    .O(net_14074)
  );
  ClkMux inmux_2_23_5_14097 (
    .I(net_5),
    .O(net_14097)
  );
  SRMux inmux_2_23_9_14098 (
    .I(net_9),
    .O(net_14098)
  );
  InMux inmux_2_2_11435_11499 (
    .I(net_11435),
    .O(net_11499)
  );
  InMux inmux_2_2_11435_11509 (
    .I(net_11435),
    .O(net_11509)
  );
  InMux inmux_2_2_11436_11498 (
    .I(net_11436),
    .O(net_11498)
  );
  InMux inmux_2_2_11436_11505 (
    .I(net_11436),
    .O(net_11505)
  );
  InMux inmux_2_2_11437_11506 (
    .I(net_11437),
    .O(net_11506)
  );
  InMux inmux_2_2_11438_11476 (
    .I(net_11438),
    .O(net_11476)
  );
  InMux inmux_2_2_11439_11492 (
    .I(net_11439),
    .O(net_11492)
  );
  InMux inmux_2_2_11440_11474 (
    .I(net_11440),
    .O(net_11474)
  );
  InMux inmux_2_2_11440_11503 (
    .I(net_11440),
    .O(net_11503)
  );
  InMux inmux_2_2_11440_11510 (
    .I(net_11440),
    .O(net_11510)
  );
  InMux inmux_2_2_11442_11511 (
    .I(net_11442),
    .O(net_11511)
  );
  InMux inmux_2_2_11444_11475 (
    .I(net_11444),
    .O(net_11475)
  );
  InMux inmux_2_2_11445_11486 (
    .I(net_11445),
    .O(net_11486)
  );
  InMux inmux_2_2_11446_11497 (
    .I(net_11446),
    .O(net_11497)
  );
  InMux inmux_2_2_11447_11479 (
    .I(net_11447),
    .O(net_11479)
  );
  InMux inmux_2_2_11448_11487 (
    .I(net_11448),
    .O(net_11487)
  );
  InMux inmux_2_2_11449_11469 (
    .I(net_11449),
    .O(net_11469)
  );
  InMux inmux_2_2_11451_11482 (
    .I(net_11451),
    .O(net_11482)
  );
  InMux inmux_2_2_11452_11488 (
    .I(net_11452),
    .O(net_11488)
  );
  InMux inmux_2_2_11454_11500 (
    .I(net_11454),
    .O(net_11500)
  );
  InMux inmux_2_2_11455_11485 (
    .I(net_11455),
    .O(net_11485)
  );
  InMux inmux_2_2_11462_11480 (
    .I(net_11462),
    .O(net_11480)
  );
  InMux inmux_2_2_11465_11481 (
    .I(net_11465),
    .O(net_11481)
  );
  ClkMux inmux_2_2_5_11514 (
    .I(net_5),
    .O(net_11514)
  );
  SRMux inmux_2_2_9_11515 (
    .I(net_9),
    .O(net_11515)
  );
  InMux inmux_2_3_11558_11603 (
    .I(net_11558),
    .O(net_11603)
  );
  InMux inmux_2_3_11560_11598 (
    .I(net_11560),
    .O(net_11598)
  );
  InMux inmux_2_3_11560_11627 (
    .I(net_11560),
    .O(net_11627)
  );
  InMux inmux_2_3_11561_11623 (
    .I(net_11561),
    .O(net_11623)
  );
  InMux inmux_2_3_11561_11633 (
    .I(net_11561),
    .O(net_11633)
  );
  InMux inmux_2_3_11562_11593 (
    .I(net_11562),
    .O(net_11593)
  );
  InMux inmux_2_3_11563_11611 (
    .I(net_11563),
    .O(net_11611)
  );
  InMux inmux_2_3_11564_11615 (
    .I(net_11564),
    .O(net_11615)
  );
  InMux inmux_2_3_11565_11620 (
    .I(net_11565),
    .O(net_11620)
  );
  InMux inmux_2_3_11565_11634 (
    .I(net_11565),
    .O(net_11634)
  );
  InMux inmux_2_3_11567_11591 (
    .I(net_11567),
    .O(net_11591)
  );
  InMux inmux_2_3_11569_11622 (
    .I(net_11569),
    .O(net_11622)
  );
  InMux inmux_2_3_11569_11632 (
    .I(net_11569),
    .O(net_11632)
  );
  InMux inmux_2_3_11570_11621 (
    .I(net_11570),
    .O(net_11621)
  );
  InMux inmux_2_3_11570_11635 (
    .I(net_11570),
    .O(net_11635)
  );
  InMux inmux_2_3_11572_11614 (
    .I(net_11572),
    .O(net_11614)
  );
  InMux inmux_2_3_11573_11597 (
    .I(net_11573),
    .O(net_11597)
  );
  InMux inmux_2_3_11573_11628 (
    .I(net_11573),
    .O(net_11628)
  );
  InMux inmux_2_3_11575_11616 (
    .I(net_11575),
    .O(net_11616)
  );
  InMux inmux_2_3_11585_11596 (
    .I(net_11585),
    .O(net_11596)
  );
  InMux inmux_2_3_11585_11629 (
    .I(net_11585),
    .O(net_11629)
  );
  InMux inmux_2_3_11586_11590 (
    .I(net_11586),
    .O(net_11590)
  );
  InMux inmux_2_3_11588_11626 (
    .I(net_11588),
    .O(net_11626)
  );
  ClkMux inmux_2_3_5_11637 (
    .I(net_5),
    .O(net_11637)
  );
  SRMux inmux_2_3_9_11638 (
    .I(net_9),
    .O(net_11638)
  );
  InMux inmux_2_4_11680_11713 (
    .I(net_11680),
    .O(net_11713)
  );
  InMux inmux_2_4_11682_11737 (
    .I(net_11682),
    .O(net_11737)
  );
  InMux inmux_2_4_11683_11731 (
    .I(net_11683),
    .O(net_11731)
  );
  InMux inmux_2_4_11683_11740 (
    .I(net_11683),
    .O(net_11740)
  );
  InMux inmux_2_4_11684_11722 (
    .I(net_11684),
    .O(net_11722)
  );
  InMux inmux_2_4_11684_11739 (
    .I(net_11684),
    .O(net_11739)
  );
  InMux inmux_2_4_11686_11732 (
    .I(net_11686),
    .O(net_11732)
  );
  InMux inmux_2_4_11690_11738 (
    .I(net_11690),
    .O(net_11738)
  );
  InMux inmux_2_4_11692_11716 (
    .I(net_11692),
    .O(net_11716)
  );
  InMux inmux_2_4_11693_11751 (
    .I(net_11693),
    .O(net_11751)
  );
  InMux inmux_2_4_11695_11756 (
    .I(net_11695),
    .O(net_11756)
  );
  InMux inmux_2_4_11696_11758 (
    .I(net_11696),
    .O(net_11758)
  );
  InMux inmux_2_4_11699_11733 (
    .I(net_11699),
    .O(net_11733)
  );
  InMux inmux_2_4_11702_11734 (
    .I(net_11702),
    .O(net_11734)
  );
  InMux inmux_2_4_11702_11749 (
    .I(net_11702),
    .O(net_11749)
  );
  InMux inmux_2_4_11704_11714 (
    .I(net_11704),
    .O(net_11714)
  );
  InMux inmux_2_4_11704_11719 (
    .I(net_11704),
    .O(net_11719)
  );
  InMux inmux_2_4_11704_11750 (
    .I(net_11704),
    .O(net_11750)
  );
  InMux inmux_2_4_11706_11745 (
    .I(net_11706),
    .O(net_11745)
  );
  InMux inmux_2_4_11707_11715 (
    .I(net_11707),
    .O(net_11715)
  );
  InMux inmux_2_4_11708_11728 (
    .I(net_11708),
    .O(net_11728)
  );
  InMux inmux_2_4_11709_11720 (
    .I(net_11709),
    .O(net_11720)
  );
  InMux inmux_2_4_11710_11755 (
    .I(net_11710),
    .O(net_11755)
  );
  ClkMux inmux_2_4_5_11760 (
    .I(net_5),
    .O(net_11760)
  );
  SRMux inmux_2_4_9_11761 (
    .I(net_9),
    .O(net_11761)
  );
  InMux inmux_2_5_11809_11855 (
    .I(net_11809),
    .O(net_11855)
  );
  InMux inmux_2_5_11816_11862 (
    .I(net_11816),
    .O(net_11862)
  );
  InMux inmux_2_5_11819_11848 (
    .I(net_11819),
    .O(net_11848)
  );
  InMux inmux_2_5_11821_11850 (
    .I(net_11821),
    .O(net_11850)
  );
  InMux inmux_2_5_11825_11838 (
    .I(net_11825),
    .O(net_11838)
  );
  InMux inmux_2_5_11829_11875 (
    .I(net_11829),
    .O(net_11875)
  );
  InMux inmux_2_5_11831_11878 (
    .I(net_11831),
    .O(net_11878)
  );
  InMux inmux_2_5_11833_11851 (
    .I(net_11833),
    .O(net_11851)
  );
  ClkMux inmux_2_5_5_11883 (
    .I(net_5),
    .O(net_11883)
  );
  SRMux inmux_2_5_9_11884 (
    .I(net_9),
    .O(net_11884)
  );
  InMux inmux_2_6_11930_11973 (
    .I(net_11930),
    .O(net_11973)
  );
  InMux inmux_2_6_11941_11995 (
    .I(net_11941),
    .O(net_11995)
  );
  InMux inmux_2_6_11943_11979 (
    .I(net_11943),
    .O(net_11979)
  );
  InMux inmux_2_6_11950_11967 (
    .I(net_11950),
    .O(net_11967)
  );
  InMux inmux_2_6_11954_11962 (
    .I(net_11954),
    .O(net_11962)
  );
  InMux inmux_2_6_11956_11991 (
    .I(net_11956),
    .O(net_11991)
  );
  InMux inmux_2_6_11957_11983 (
    .I(net_11957),
    .O(net_11983)
  );
  ClkMux inmux_2_6_5_12006 (
    .I(net_5),
    .O(net_12006)
  );
  SRMux inmux_2_6_9_12007 (
    .I(net_9),
    .O(net_12007)
  );
  InMux inmux_2_7_12050_12088 (
    .I(net_12050),
    .O(net_12088)
  );
  InMux inmux_2_7_12053_12089 (
    .I(net_12053),
    .O(net_12089)
  );
  InMux inmux_2_7_12054_12100 (
    .I(net_12054),
    .O(net_12100)
  );
  InMux inmux_2_7_12056_12083 (
    .I(net_12056),
    .O(net_12083)
  );
  InMux inmux_2_7_12065_12106 (
    .I(net_12065),
    .O(net_12106)
  );
  InMux inmux_2_7_12067_12091 (
    .I(net_12067),
    .O(net_12091)
  );
  InMux inmux_2_7_12071_12120 (
    .I(net_12071),
    .O(net_12120)
  );
  InMux inmux_2_7_12073_12090 (
    .I(net_12073),
    .O(net_12090)
  );
  InMux inmux_2_7_12077_12124 (
    .I(net_12077),
    .O(net_12124)
  );
  ClkMux inmux_2_7_5_12129 (
    .I(net_5),
    .O(net_12129)
  );
  CEMux inmux_2_7_8_12128 (
    .I(net_8),
    .O(net_12128)
  );
  InMux inmux_2_8_12172_12231 (
    .I(net_12172),
    .O(net_12231)
  );
  CEMux inmux_2_8_12174_12251 (
    .I(net_12174),
    .O(net_12251)
  );
  InMux inmux_2_8_12175_12211 (
    .I(net_12175),
    .O(net_12211)
  );
  InMux inmux_2_8_12176_12226 (
    .I(net_12176),
    .O(net_12226)
  );
  InMux inmux_2_8_12177_12230 (
    .I(net_12177),
    .O(net_12230)
  );
  InMux inmux_2_8_12178_12238 (
    .I(net_12178),
    .O(net_12238)
  );
  InMux inmux_2_8_12179_12213 (
    .I(net_12179),
    .O(net_12213)
  );
  InMux inmux_2_8_12180_12206 (
    .I(net_12180),
    .O(net_12206)
  );
  InMux inmux_2_8_12180_12223 (
    .I(net_12180),
    .O(net_12223)
  );
  InMux inmux_2_8_12181_12205 (
    .I(net_12181),
    .O(net_12205)
  );
  InMux inmux_2_8_12181_12212 (
    .I(net_12181),
    .O(net_12212)
  );
  InMux inmux_2_8_12182_12225 (
    .I(net_12182),
    .O(net_12225)
  );
  InMux inmux_2_8_12182_12232 (
    .I(net_12182),
    .O(net_12232)
  );
  InMux inmux_2_8_12183_12214 (
    .I(net_12183),
    .O(net_12214)
  );
  InMux inmux_2_8_12184_12220 (
    .I(net_12184),
    .O(net_12220)
  );
  InMux inmux_2_8_12186_12208 (
    .I(net_12186),
    .O(net_12208)
  );
  InMux inmux_2_8_12187_12229 (
    .I(net_12187),
    .O(net_12229)
  );
  InMux inmux_2_8_12190_12207 (
    .I(net_12190),
    .O(net_12207)
  );
  InMux inmux_2_8_12193_12249 (
    .I(net_12193),
    .O(net_12249)
  );
  InMux inmux_2_8_12194_12224 (
    .I(net_12194),
    .O(net_12224)
  );
  InMux inmux_2_8_12201_12241 (
    .I(net_12201),
    .O(net_12241)
  );
  ClkMux inmux_2_8_5_12252 (
    .I(net_5),
    .O(net_12252)
  );
  InMux inmux_2_9_12295_12364 (
    .I(net_12295),
    .O(net_12364)
  );
  InMux inmux_2_9_12297_12328 (
    .I(net_12297),
    .O(net_12328)
  );
  InMux inmux_2_9_12299_12373 (
    .I(net_12299),
    .O(net_12373)
  );
  InMux inmux_2_9_12300_12358 (
    .I(net_12300),
    .O(net_12358)
  );
  InMux inmux_2_9_12302_12346 (
    .I(net_12302),
    .O(net_12346)
  );
  InMux inmux_2_9_12308_12352 (
    .I(net_12308),
    .O(net_12352)
  );
  InMux inmux_2_9_12312_12334 (
    .I(net_12312),
    .O(net_12334)
  );
  InMux inmux_2_9_12319_12343 (
    .I(net_12319),
    .O(net_12343)
  );
  ClkMux inmux_2_9_5_12375 (
    .I(net_5),
    .O(net_12375)
  );
  SRMux inmux_2_9_9_12376 (
    .I(net_9),
    .O(net_12376)
  );
  InMux inmux_3_10_16253_16315 (
    .I(net_16253),
    .O(net_16315)
  );
  InMux inmux_3_10_16254_16300 (
    .I(net_16254),
    .O(net_16300)
  );
  InMux inmux_3_10_16260_16291 (
    .I(net_16260),
    .O(net_16291)
  );
  InMux inmux_3_10_16261_16309 (
    .I(net_16261),
    .O(net_16309)
  );
  InMux inmux_3_10_16268_16326 (
    .I(net_16268),
    .O(net_16326)
  );
  InMux inmux_3_10_16273_16283 (
    .I(net_16273),
    .O(net_16283)
  );
  InMux inmux_3_10_16276_16320 (
    .I(net_16276),
    .O(net_16320)
  );
  InMux inmux_3_10_16278_16296 (
    .I(net_16278),
    .O(net_16296)
  );
  ClkMux inmux_3_10_5_16329 (
    .I(net_5),
    .O(net_16329)
  );
  SRMux inmux_3_10_9_16330 (
    .I(net_9),
    .O(net_16330)
  );
  InMux inmux_3_11_16375_16425 (
    .I(net_16375),
    .O(net_16425)
  );
  InMux inmux_3_11_16383_16414 (
    .I(net_16383),
    .O(net_16414)
  );
  InMux inmux_3_11_16385_16431 (
    .I(net_16385),
    .O(net_16431)
  );
  InMux inmux_3_11_16386_16406 (
    .I(net_16386),
    .O(net_16406)
  );
  InMux inmux_3_11_16387_16443 (
    .I(net_16387),
    .O(net_16443)
  );
  InMux inmux_3_11_16388_16419 (
    .I(net_16388),
    .O(net_16419)
  );
  InMux inmux_3_11_16390_16450 (
    .I(net_16390),
    .O(net_16450)
  );
  InMux inmux_3_11_16394_16436 (
    .I(net_16394),
    .O(net_16436)
  );
  ClkMux inmux_3_11_5_16452 (
    .I(net_5),
    .O(net_16452)
  );
  SRMux inmux_3_11_9_16453 (
    .I(net_9),
    .O(net_16453)
  );
  InMux inmux_3_12_16498_16536 (
    .I(net_16498),
    .O(net_16536)
  );
  InMux inmux_3_12_16499_16547 (
    .I(net_16499),
    .O(net_16547)
  );
  InMux inmux_3_12_16500_16529 (
    .I(net_16500),
    .O(net_16529)
  );
  InMux inmux_3_12_16504_16542 (
    .I(net_16504),
    .O(net_16542)
  );
  InMux inmux_3_12_16507_16560 (
    .I(net_16507),
    .O(net_16560)
  );
  InMux inmux_3_12_16508_16559 (
    .I(net_16508),
    .O(net_16559)
  );
  InMux inmux_3_12_16510_16535 (
    .I(net_16510),
    .O(net_16535)
  );
  InMux inmux_3_12_16513_16566 (
    .I(net_16513),
    .O(net_16566)
  );
  InMux inmux_3_12_16514_16553 (
    .I(net_16514),
    .O(net_16553)
  );
  InMux inmux_3_12_16515_16554 (
    .I(net_16515),
    .O(net_16554)
  );
  InMux inmux_3_12_16517_16530 (
    .I(net_16517),
    .O(net_16530)
  );
  InMux inmux_3_12_16518_16565 (
    .I(net_16518),
    .O(net_16565)
  );
  InMux inmux_3_12_16523_16541 (
    .I(net_16523),
    .O(net_16541)
  );
  InMux inmux_3_12_16525_16548 (
    .I(net_16525),
    .O(net_16548)
  );
  InMux inmux_3_12_16527_16537 (
    .I(net_16527),
    .O(net_16537)
  );
  InMux inmux_3_12_16533_16543 (
    .I(net_16533),
    .O(net_16543)
  );
  InMux inmux_3_12_16539_16549 (
    .I(net_16539),
    .O(net_16549)
  );
  InMux inmux_3_12_16545_16555 (
    .I(net_16545),
    .O(net_16555)
  );
  InMux inmux_3_12_16551_16561 (
    .I(net_16551),
    .O(net_16561)
  );
  InMux inmux_3_12_16557_16567 (
    .I(net_16557),
    .O(net_16567)
  );
  InMux inmux_3_12_16563_16573 (
    .I(net_16563),
    .O(net_16573)
  );
  InMux inmux_3_13_16623_16652 (
    .I(net_16623),
    .O(net_16652)
  );
  InMux inmux_3_13_16625_16671 (
    .I(net_16625),
    .O(net_16671)
  );
  InMux inmux_3_13_16633_16653 (
    .I(net_16633),
    .O(net_16653)
  );
  InMux inmux_3_13_16634_16677 (
    .I(net_16634),
    .O(net_16677)
  );
  InMux inmux_3_13_16636_16670 (
    .I(net_16636),
    .O(net_16670)
  );
  InMux inmux_3_13_16637_16676 (
    .I(net_16637),
    .O(net_16676)
  );
  InMux inmux_3_13_16638_16682 (
    .I(net_16638),
    .O(net_16682)
  );
  InMux inmux_3_13_16639_16688 (
    .I(net_16639),
    .O(net_16688)
  );
  InMux inmux_3_13_16640_16694 (
    .I(net_16640),
    .O(net_16694)
  );
  InMux inmux_3_13_16642_16659 (
    .I(net_16642),
    .O(net_16659)
  );
  InMux inmux_3_13_16643_16665 (
    .I(net_16643),
    .O(net_16665)
  );
  InMux inmux_3_13_16644_16683 (
    .I(net_16644),
    .O(net_16683)
  );
  InMux inmux_3_13_16645_16658 (
    .I(net_16645),
    .O(net_16658)
  );
  InMux inmux_3_13_16646_16664 (
    .I(net_16646),
    .O(net_16664)
  );
  InMux inmux_3_13_16647_16689 (
    .I(net_16647),
    .O(net_16689)
  );
  InMux inmux_3_13_16648_16695 (
    .I(net_16648),
    .O(net_16695)
  );
  InMux inmux_3_13_16650_16660 (
    .I(net_16650),
    .O(net_16660)
  );
  InMux inmux_3_13_16656_16666 (
    .I(net_16656),
    .O(net_16666)
  );
  InMux inmux_3_13_16662_16672 (
    .I(net_16662),
    .O(net_16672)
  );
  InMux inmux_3_13_16668_16678 (
    .I(net_16668),
    .O(net_16678)
  );
  InMux inmux_3_13_16674_16684 (
    .I(net_16674),
    .O(net_16684)
  );
  InMux inmux_3_13_16680_16690 (
    .I(net_16680),
    .O(net_16690)
  );
  InMux inmux_3_13_16686_16696 (
    .I(net_16686),
    .O(net_16696)
  );
  ClkMux inmux_3_13_5_16698 (
    .I(net_5),
    .O(net_16698)
  );
  SRMux inmux_3_13_9_16699 (
    .I(net_9),
    .O(net_16699)
  );
  InMux inmux_3_14_16736_16777 (
    .I(net_16736),
    .O(net_16777)
  );
  InMux inmux_3_14_16742_16804 (
    .I(net_16742),
    .O(net_16804)
  );
  InMux inmux_3_14_16748_16775 (
    .I(net_16748),
    .O(net_16775)
  );
  InMux inmux_3_14_16748_16782 (
    .I(net_16748),
    .O(net_16782)
  );
  InMux inmux_3_14_16756_16776 (
    .I(net_16756),
    .O(net_16776)
  );
  InMux inmux_3_14_16757_16817 (
    .I(net_16757),
    .O(net_16817)
  );
  InMux inmux_3_14_16758_16799 (
    .I(net_16758),
    .O(net_16799)
  );
  InMux inmux_3_14_16761_16807 (
    .I(net_16761),
    .O(net_16807)
  );
  InMux inmux_3_14_16762_16787 (
    .I(net_16762),
    .O(net_16787)
  );
  InMux inmux_3_14_16765_16780 (
    .I(net_16765),
    .O(net_16780)
  );
  InMux inmux_3_14_16767_16794 (
    .I(net_16767),
    .O(net_16794)
  );
  InMux inmux_3_14_16768_16805 (
    .I(net_16768),
    .O(net_16805)
  );
  InMux inmux_3_14_16770_16812 (
    .I(net_16770),
    .O(net_16812)
  );
  InMux inmux_3_14_16773_16783 (
    .I(net_16773),
    .O(net_16783)
  );
  ClkMux inmux_3_14_5_16821 (
    .I(net_5),
    .O(net_16821)
  );
  SRMux inmux_3_14_9_16822 (
    .I(net_9),
    .O(net_16822)
  );
  InMux inmux_3_15_16864_16928 (
    .I(net_16864),
    .O(net_16928)
  );
  InMux inmux_3_15_16866_16899 (
    .I(net_16866),
    .O(net_16899)
  );
  InMux inmux_3_15_16867_16898 (
    .I(net_16867),
    .O(net_16898)
  );
  InMux inmux_3_15_16868_16916 (
    .I(net_16868),
    .O(net_16916)
  );
  InMux inmux_3_15_16869_16929 (
    .I(net_16869),
    .O(net_16929)
  );
  InMux inmux_3_15_16873_16935 (
    .I(net_16873),
    .O(net_16935)
  );
  InMux inmux_3_15_16878_16922 (
    .I(net_16878),
    .O(net_16922)
  );
  InMux inmux_3_15_16883_16917 (
    .I(net_16883),
    .O(net_16917)
  );
  InMux inmux_3_15_16884_16923 (
    .I(net_16884),
    .O(net_16923)
  );
  InMux inmux_3_15_16886_16911 (
    .I(net_16886),
    .O(net_16911)
  );
  InMux inmux_3_15_16890_16910 (
    .I(net_16890),
    .O(net_16910)
  );
  InMux inmux_3_15_16892_16905 (
    .I(net_16892),
    .O(net_16905)
  );
  InMux inmux_3_15_16893_16904 (
    .I(net_16893),
    .O(net_16904)
  );
  InMux inmux_3_15_16894_16934 (
    .I(net_16894),
    .O(net_16934)
  );
  InMux inmux_3_15_16896_16906 (
    .I(net_16896),
    .O(net_16906)
  );
  InMux inmux_3_15_16902_16912 (
    .I(net_16902),
    .O(net_16912)
  );
  InMux inmux_3_15_16908_16918 (
    .I(net_16908),
    .O(net_16918)
  );
  InMux inmux_3_15_16914_16924 (
    .I(net_16914),
    .O(net_16924)
  );
  InMux inmux_3_15_16920_16930 (
    .I(net_16920),
    .O(net_16930)
  );
  InMux inmux_3_15_16926_16936 (
    .I(net_16926),
    .O(net_16936)
  );
  InMux inmux_3_15_16932_16942 (
    .I(net_16932),
    .O(net_16942)
  );
  InMux inmux_3_16_16989_17041 (
    .I(net_16989),
    .O(net_17041)
  );
  InMux inmux_3_16_16990_17057 (
    .I(net_16990),
    .O(net_17057)
  );
  InMux inmux_3_16_16992_17023 (
    .I(net_16992),
    .O(net_17023)
  );
  InMux inmux_3_16_16998_17051 (
    .I(net_16998),
    .O(net_17051)
  );
  InMux inmux_3_16_16999_17045 (
    .I(net_16999),
    .O(net_17045)
  );
  InMux inmux_3_16_17001_17033 (
    .I(net_17001),
    .O(net_17033)
  );
  InMux inmux_3_16_17004_17062 (
    .I(net_17004),
    .O(net_17062)
  );
  InMux inmux_3_16_17016_17029 (
    .I(net_17016),
    .O(net_17029)
  );
  ClkMux inmux_3_16_5_17067 (
    .I(net_5),
    .O(net_17067)
  );
  SRMux inmux_3_16_9_17068 (
    .I(net_9),
    .O(net_17068)
  );
  InMux inmux_3_17_17114_17143 (
    .I(net_17114),
    .O(net_17143)
  );
  InMux inmux_3_17_17115_17173 (
    .I(net_17115),
    .O(net_17173)
  );
  InMux inmux_3_17_17121_17169 (
    .I(net_17121),
    .O(net_17169)
  );
  InMux inmux_3_17_17126_17164 (
    .I(net_17126),
    .O(net_17164)
  );
  InMux inmux_3_17_17127_17158 (
    .I(net_17127),
    .O(net_17158)
  );
  InMux inmux_3_17_17132_17179 (
    .I(net_17132),
    .O(net_17179)
  );
  InMux inmux_3_17_17133_17185 (
    .I(net_17133),
    .O(net_17185)
  );
  ClkMux inmux_3_17_5_17190 (
    .I(net_5),
    .O(net_17190)
  );
  SRMux inmux_3_17_9_17191 (
    .I(net_9),
    .O(net_17191)
  );
  InMux inmux_3_18_17233_17268 (
    .I(net_17233),
    .O(net_17268)
  );
  InMux inmux_3_18_17234_17296 (
    .I(net_17234),
    .O(net_17296)
  );
  InMux inmux_3_18_17234_17303 (
    .I(net_17234),
    .O(net_17303)
  );
  InMux inmux_3_18_17237_17304 (
    .I(net_17237),
    .O(net_17304)
  );
  InMux inmux_3_18_17238_17291 (
    .I(net_17238),
    .O(net_17291)
  );
  InMux inmux_3_18_17241_17298 (
    .I(net_17241),
    .O(net_17298)
  );
  InMux inmux_3_18_17242_17302 (
    .I(net_17242),
    .O(net_17302)
  );
  InMux inmux_3_18_17243_17305 (
    .I(net_17243),
    .O(net_17305)
  );
  CEMux inmux_3_18_17244_17312 (
    .I(net_17244),
    .O(net_17312)
  );
  InMux inmux_3_18_17245_17267 (
    .I(net_17245),
    .O(net_17267)
  );
  InMux inmux_3_18_17246_17299 (
    .I(net_17246),
    .O(net_17299)
  );
  InMux inmux_3_18_17248_17297 (
    .I(net_17248),
    .O(net_17297)
  );
  InMux inmux_3_18_17249_17266 (
    .I(net_17249),
    .O(net_17266)
  );
  InMux inmux_3_18_17253_17309 (
    .I(net_17253),
    .O(net_17309)
  );
  InMux inmux_3_18_17259_17269 (
    .I(net_17259),
    .O(net_17269)
  );
  ClkMux inmux_3_18_5_17313 (
    .I(net_5),
    .O(net_17313)
  );
  SRMux inmux_3_18_9_17314 (
    .I(net_9),
    .O(net_17314)
  );
  InMux inmux_3_19_17364_17402 (
    .I(net_17364),
    .O(net_17402)
  );
  InMux inmux_3_19_17373_17421 (
    .I(net_17373),
    .O(net_17421)
  );
  ClkMux inmux_3_19_5_17436 (
    .I(net_5),
    .O(net_17436)
  );
  SRMux inmux_3_19_9_17437 (
    .I(net_9),
    .O(net_17437)
  );
  InMux inmux_3_1_15103_15136 (
    .I(net_15103),
    .O(net_15136)
  );
  CEMux inmux_3_1_15104_15181 (
    .I(net_15104),
    .O(net_15181)
  );
  InMux inmux_3_1_15106_15149 (
    .I(net_15106),
    .O(net_15149)
  );
  InMux inmux_3_1_15110_15143 (
    .I(net_15110),
    .O(net_15143)
  );
  InMux inmux_3_1_15115_15156 (
    .I(net_15115),
    .O(net_15156)
  );
  InMux inmux_3_1_15118_15142 (
    .I(net_15118),
    .O(net_15142)
  );
  InMux inmux_3_1_15119_15138 (
    .I(net_15119),
    .O(net_15138)
  );
  InMux inmux_3_1_15119_15155 (
    .I(net_15119),
    .O(net_15155)
  );
  InMux inmux_3_1_15120_15180 (
    .I(net_15120),
    .O(net_15180)
  );
  InMux inmux_3_1_15121_15141 (
    .I(net_15121),
    .O(net_15141)
  );
  InMux inmux_3_1_15121_15150 (
    .I(net_15121),
    .O(net_15150)
  );
  InMux inmux_3_1_15121_15153 (
    .I(net_15121),
    .O(net_15153)
  );
  InMux inmux_3_1_15121_15177 (
    .I(net_15121),
    .O(net_15177)
  );
  InMux inmux_3_1_15122_15137 (
    .I(net_15122),
    .O(net_15137)
  );
  InMux inmux_3_1_15124_15135 (
    .I(net_15124),
    .O(net_15135)
  );
  InMux inmux_3_1_15126_15179 (
    .I(net_15126),
    .O(net_15179)
  );
  InMux inmux_3_1_15127_15147 (
    .I(net_15127),
    .O(net_15147)
  );
  InMux inmux_3_1_15127_15178 (
    .I(net_15127),
    .O(net_15178)
  );
  InMux inmux_3_1_15129_15173 (
    .I(net_15129),
    .O(net_15173)
  );
  InMux inmux_3_1_15131_15171 (
    .I(net_15131),
    .O(net_15171)
  );
  InMux inmux_3_1_15132_15148 (
    .I(net_15132),
    .O(net_15148)
  );
  InMux inmux_3_1_15133_15154 (
    .I(net_15133),
    .O(net_15154)
  );
  ClkMux inmux_3_1_5_15182 (
    .I(net_5),
    .O(net_15182)
  );
  SRMux inmux_3_1_9_15183 (
    .I(net_9),
    .O(net_15183)
  );
  InMux inmux_3_20_17504_17521 (
    .I(net_17504),
    .O(net_17521)
  );
  ClkMux inmux_3_20_5_17559 (
    .I(net_5),
    .O(net_17559)
  );
  SRMux inmux_3_20_9_17560 (
    .I(net_9),
    .O(net_17560)
  );
  InMux inmux_3_21_17613_17666 (
    .I(net_17613),
    .O(net_17666)
  );
  InMux inmux_3_21_17620_17671 (
    .I(net_17620),
    .O(net_17671)
  );
  ClkMux inmux_3_21_5_17682 (
    .I(net_5),
    .O(net_17682)
  );
  SRMux inmux_3_21_9_17683 (
    .I(net_9),
    .O(net_17683)
  );
  InMux inmux_3_22_17745_17777 (
    .I(net_17745),
    .O(net_17777)
  );
  ClkMux inmux_3_22_5_17805 (
    .I(net_5),
    .O(net_17805)
  );
  SRMux inmux_3_22_9_17806 (
    .I(net_9),
    .O(net_17806)
  );
  InMux inmux_3_2_15265_15317 (
    .I(net_15265),
    .O(net_15317)
  );
  InMux inmux_3_2_15268_15311 (
    .I(net_15268),
    .O(net_15311)
  );
  InMux inmux_3_2_15268_15323 (
    .I(net_15268),
    .O(net_15323)
  );
  InMux inmux_3_2_15268_15342 (
    .I(net_15268),
    .O(net_15342)
  );
  InMux inmux_3_2_15269_15298 (
    .I(net_15269),
    .O(net_15298)
  );
  InMux inmux_3_2_15270_15301 (
    .I(net_15270),
    .O(net_15301)
  );
  InMux inmux_3_2_15270_15306 (
    .I(net_15270),
    .O(net_15306)
  );
  InMux inmux_3_2_15270_15328 (
    .I(net_15270),
    .O(net_15328)
  );
  InMux inmux_3_2_15273_15335 (
    .I(net_15273),
    .O(net_15335)
  );
  InMux inmux_3_2_15274_15312 (
    .I(net_15274),
    .O(net_15312)
  );
  InMux inmux_3_2_15279_15316 (
    .I(net_15279),
    .O(net_15316)
  );
  InMux inmux_3_2_15280_15322 (
    .I(net_15280),
    .O(net_15322)
  );
  InMux inmux_3_2_15282_15299 (
    .I(net_15282),
    .O(net_15299)
  );
  CEMux inmux_3_2_15283_15344 (
    .I(net_15283),
    .O(net_15344)
  );
  InMux inmux_3_2_15284_15337 (
    .I(net_15284),
    .O(net_15337)
  );
  InMux inmux_3_2_15285_15305 (
    .I(net_15285),
    .O(net_15305)
  );
  InMux inmux_3_2_15286_15330 (
    .I(net_15286),
    .O(net_15330)
  );
  InMux inmux_3_2_15289_15325 (
    .I(net_15289),
    .O(net_15325)
  );
  InMux inmux_3_2_15290_15300 (
    .I(net_15290),
    .O(net_15300)
  );
  InMux inmux_3_2_15290_15307 (
    .I(net_15290),
    .O(net_15307)
  );
  InMux inmux_3_2_15290_15319 (
    .I(net_15290),
    .O(net_15319)
  );
  InMux inmux_3_2_15290_15329 (
    .I(net_15290),
    .O(net_15329)
  );
  InMux inmux_3_2_15291_15304 (
    .I(net_15291),
    .O(net_15304)
  );
  InMux inmux_3_2_15292_15343 (
    .I(net_15292),
    .O(net_15343)
  );
  InMux inmux_3_2_15293_15313 (
    .I(net_15293),
    .O(net_15313)
  );
  InMux inmux_3_2_15294_15341 (
    .I(net_15294),
    .O(net_15341)
  );
  InMux inmux_3_2_15295_15318 (
    .I(net_15295),
    .O(net_15318)
  );
  InMux inmux_3_2_15296_15331 (
    .I(net_15296),
    .O(net_15331)
  );
  ClkMux inmux_3_2_5_15345 (
    .I(net_5),
    .O(net_15345)
  );
  SRMux inmux_3_2_9_15346 (
    .I(net_9),
    .O(net_15346)
  );
  InMux inmux_3_3_15390_15442 (
    .I(net_15390),
    .O(net_15442)
  );
  InMux inmux_3_3_15390_15466 (
    .I(net_15390),
    .O(net_15466)
  );
  CEMux inmux_3_3_15390_15467 (
    .I(net_15390),
    .O(net_15467)
  );
  InMux inmux_3_3_15391_15458 (
    .I(net_15391),
    .O(net_15458)
  );
  InMux inmux_3_3_15392_15445 (
    .I(net_15392),
    .O(net_15445)
  );
  InMux inmux_3_3_15394_15423 (
    .I(net_15394),
    .O(net_15423)
  );
  InMux inmux_3_3_15395_15448 (
    .I(net_15395),
    .O(net_15448)
  );
  InMux inmux_3_3_15397_15433 (
    .I(net_15397),
    .O(net_15433)
  );
  InMux inmux_3_3_15398_15427 (
    .I(net_15398),
    .O(net_15427)
  );
  InMux inmux_3_3_15398_15460 (
    .I(net_15398),
    .O(net_15460)
  );
  InMux inmux_3_3_15399_15454 (
    .I(net_15399),
    .O(net_15454)
  );
  InMux inmux_3_3_15400_15439 (
    .I(net_15400),
    .O(net_15439)
  );
  InMux inmux_3_3_15402_15434 (
    .I(net_15402),
    .O(net_15434)
  );
  InMux inmux_3_3_15404_15459 (
    .I(net_15404),
    .O(net_15459)
  );
  InMux inmux_3_3_15406_15452 (
    .I(net_15406),
    .O(net_15452)
  );
  InMux inmux_3_3_15407_15422 (
    .I(net_15407),
    .O(net_15422)
  );
  InMux inmux_3_3_15407_15429 (
    .I(net_15407),
    .O(net_15429)
  );
  InMux inmux_3_3_15407_15453 (
    .I(net_15407),
    .O(net_15453)
  );
  InMux inmux_3_3_15408_15421 (
    .I(net_15408),
    .O(net_15421)
  );
  InMux inmux_3_3_15409_15441 (
    .I(net_15409),
    .O(net_15441)
  );
  InMux inmux_3_3_15410_15440 (
    .I(net_15410),
    .O(net_15440)
  );
  InMux inmux_3_3_15410_15447 (
    .I(net_15410),
    .O(net_15447)
  );
  InMux inmux_3_3_15412_15465 (
    .I(net_15412),
    .O(net_15465)
  );
  InMux inmux_3_3_15414_15424 (
    .I(net_15414),
    .O(net_15424)
  );
  InMux inmux_3_3_15414_15451 (
    .I(net_15414),
    .O(net_15451)
  );
  InMux inmux_3_3_15415_15430 (
    .I(net_15415),
    .O(net_15430)
  );
  InMux inmux_3_3_15416_15463 (
    .I(net_15416),
    .O(net_15463)
  );
  InMux inmux_3_3_15417_15428 (
    .I(net_15417),
    .O(net_15428)
  );
  InMux inmux_3_3_15417_15457 (
    .I(net_15417),
    .O(net_15457)
  );
  InMux inmux_3_3_15417_15464 (
    .I(net_15417),
    .O(net_15464)
  );
  ClkMux inmux_3_3_5_15468 (
    .I(net_5),
    .O(net_15468)
  );
  SRMux inmux_3_3_9_15469 (
    .I(net_9),
    .O(net_15469)
  );
  InMux inmux_3_4_15511_15568 (
    .I(net_15511),
    .O(net_15568)
  );
  InMux inmux_3_4_15514_15569 (
    .I(net_15514),
    .O(net_15569)
  );
  InMux inmux_3_4_15516_15547 (
    .I(net_15516),
    .O(net_15547)
  );
  InMux inmux_3_4_15518_15545 (
    .I(net_15518),
    .O(net_15545)
  );
  InMux inmux_3_4_15519_15574 (
    .I(net_15519),
    .O(net_15574)
  );
  InMux inmux_3_4_15522_15587 (
    .I(net_15522),
    .O(net_15587)
  );
  InMux inmux_3_4_15523_15564 (
    .I(net_15523),
    .O(net_15564)
  );
  InMux inmux_3_4_15524_15570 (
    .I(net_15524),
    .O(net_15570)
  );
  InMux inmux_3_4_15525_15583 (
    .I(net_15525),
    .O(net_15583)
  );
  InMux inmux_3_4_15526_15577 (
    .I(net_15526),
    .O(net_15577)
  );
  InMux inmux_3_4_15526_15589 (
    .I(net_15526),
    .O(net_15589)
  );
  InMux inmux_3_4_15527_15556 (
    .I(net_15527),
    .O(net_15556)
  );
  InMux inmux_3_4_15530_15557 (
    .I(net_15530),
    .O(net_15557)
  );
  InMux inmux_3_4_15533_15544 (
    .I(net_15533),
    .O(net_15544)
  );
  InMux inmux_3_4_15533_15575 (
    .I(net_15533),
    .O(net_15575)
  );
  InMux inmux_3_4_15536_15546 (
    .I(net_15536),
    .O(net_15546)
  );
  ClkMux inmux_3_4_5_15591 (
    .I(net_5),
    .O(net_15591)
  );
  SRMux inmux_3_4_9_15592 (
    .I(net_9),
    .O(net_15592)
  );
  InMux inmux_3_5_15638_15674 (
    .I(net_15638),
    .O(net_15674)
  );
  InMux inmux_3_5_15640_15705 (
    .I(net_15640),
    .O(net_15705)
  );
  InMux inmux_3_5_15642_15668 (
    .I(net_15642),
    .O(net_15668)
  );
  InMux inmux_3_5_15644_15709 (
    .I(net_15644),
    .O(net_15709)
  );
  InMux inmux_3_5_15648_15670 (
    .I(net_15648),
    .O(net_15670)
  );
  InMux inmux_3_5_15651_15682 (
    .I(net_15651),
    .O(net_15682)
  );
  InMux inmux_3_5_15653_15692 (
    .I(net_15653),
    .O(net_15692)
  );
  InMux inmux_3_5_15655_15694 (
    .I(net_15655),
    .O(net_15694)
  );
  InMux inmux_3_5_15660_15697 (
    .I(net_15660),
    .O(net_15697)
  );
  ClkMux inmux_3_5_5_15714 (
    .I(net_5),
    .O(net_15714)
  );
  SRMux inmux_3_5_9_15715 (
    .I(net_9),
    .O(net_15715)
  );
  InMux inmux_3_6_15761_15814 (
    .I(net_15761),
    .O(net_15814)
  );
  InMux inmux_3_6_15762_15791 (
    .I(net_15762),
    .O(net_15791)
  );
  InMux inmux_3_6_15765_15829 (
    .I(net_15765),
    .O(net_15829)
  );
  InMux inmux_3_6_15766_15797 (
    .I(net_15766),
    .O(net_15797)
  );
  InMux inmux_3_6_15767_15820 (
    .I(net_15767),
    .O(net_15820)
  );
  InMux inmux_3_6_15770_15828 (
    .I(net_15770),
    .O(net_15828)
  );
  InMux inmux_3_6_15772_15816 (
    .I(net_15772),
    .O(net_15816)
  );
  InMux inmux_3_6_15774_15817 (
    .I(net_15774),
    .O(net_15817)
  );
  CEMux inmux_3_6_15775_15836 (
    .I(net_15775),
    .O(net_15836)
  );
  InMux inmux_3_6_15776_15827 (
    .I(net_15776),
    .O(net_15827)
  );
  InMux inmux_3_6_15781_15815 (
    .I(net_15781),
    .O(net_15815)
  );
  InMux inmux_3_6_15783_15808 (
    .I(net_15783),
    .O(net_15808)
  );
  InMux inmux_3_6_15784_15835 (
    .I(net_15784),
    .O(net_15835)
  );
  ClkMux inmux_3_6_5_15837 (
    .I(net_5),
    .O(net_15837)
  );
  InMux inmux_3_7_15882_15939 (
    .I(net_15882),
    .O(net_15939)
  );
  InMux inmux_3_7_15883_15938 (
    .I(net_15883),
    .O(net_15938)
  );
  InMux inmux_3_7_15884_15944 (
    .I(net_15884),
    .O(net_15944)
  );
  InMux inmux_3_7_15885_15933 (
    .I(net_15885),
    .O(net_15933)
  );
  InMux inmux_3_7_15886_15920 (
    .I(net_15886),
    .O(net_15920)
  );
  InMux inmux_3_7_15888_15914 (
    .I(net_15888),
    .O(net_15914)
  );
  InMux inmux_3_7_15888_15957 (
    .I(net_15888),
    .O(net_15957)
  );
  InMux inmux_3_7_15889_15915 (
    .I(net_15889),
    .O(net_15915)
  );
  InMux inmux_3_7_15889_15956 (
    .I(net_15889),
    .O(net_15956)
  );
  InMux inmux_3_7_15890_15945 (
    .I(net_15890),
    .O(net_15945)
  );
  InMux inmux_3_7_15891_15927 (
    .I(net_15891),
    .O(net_15927)
  );
  InMux inmux_3_7_15892_15921 (
    .I(net_15892),
    .O(net_15921)
  );
  InMux inmux_3_7_15894_15926 (
    .I(net_15894),
    .O(net_15926)
  );
  InMux inmux_3_7_15895_15932 (
    .I(net_15895),
    .O(net_15932)
  );
  InMux inmux_3_7_15912_15922 (
    .I(net_15912),
    .O(net_15922)
  );
  InMux inmux_3_7_15918_15928 (
    .I(net_15918),
    .O(net_15928)
  );
  InMux inmux_3_7_15924_15934 (
    .I(net_15924),
    .O(net_15934)
  );
  InMux inmux_3_7_15930_15940 (
    .I(net_15930),
    .O(net_15940)
  );
  InMux inmux_3_7_15936_15946 (
    .I(net_15936),
    .O(net_15946)
  );
  InMux inmux_3_7_15942_15952 (
    .I(net_15942),
    .O(net_15952)
  );
  ClkMux inmux_3_7_5_15960 (
    .I(net_5),
    .O(net_15960)
  );
  SRMux inmux_3_7_9_15961 (
    .I(net_9),
    .O(net_15961)
  );
  CEMux inmux_3_8_12_16082 (
    .I(net_12),
    .O(net_16082)
  );
  InMux inmux_3_8_16003_16079 (
    .I(net_16003),
    .O(net_16079)
  );
  InMux inmux_3_8_16005_16038 (
    .I(net_16005),
    .O(net_16038)
  );
  InMux inmux_3_8_16013_16063 (
    .I(net_16013),
    .O(net_16063)
  );
  InMux inmux_3_8_16020_16061 (
    .I(net_16020),
    .O(net_16061)
  );
  InMux inmux_3_8_16023_16060 (
    .I(net_16023),
    .O(net_16060)
  );
  InMux inmux_3_8_16029_16051 (
    .I(net_16029),
    .O(net_16051)
  );
  ClkMux inmux_3_8_5_16083 (
    .I(net_5),
    .O(net_16083)
  );
  InMux inmux_3_9_16127_16196 (
    .I(net_16127),
    .O(net_16196)
  );
  InMux inmux_3_9_16129_16184 (
    .I(net_16129),
    .O(net_16184)
  );
  InMux inmux_3_9_16130_16190 (
    .I(net_16130),
    .O(net_16190)
  );
  InMux inmux_3_9_16132_16185 (
    .I(net_16132),
    .O(net_16185)
  );
  InMux inmux_3_9_16133_16191 (
    .I(net_16133),
    .O(net_16191)
  );
  InMux inmux_3_9_16134_16172 (
    .I(net_16134),
    .O(net_16172)
  );
  InMux inmux_3_9_16135_16161 (
    .I(net_16135),
    .O(net_16161)
  );
  InMux inmux_3_9_16138_16160 (
    .I(net_16138),
    .O(net_16160)
  );
  InMux inmux_3_9_16139_16178 (
    .I(net_16139),
    .O(net_16178)
  );
  InMux inmux_3_9_16141_16166 (
    .I(net_16141),
    .O(net_16166)
  );
  InMux inmux_3_9_16142_16197 (
    .I(net_16142),
    .O(net_16197)
  );
  InMux inmux_3_9_16149_16167 (
    .I(net_16149),
    .O(net_16167)
  );
  InMux inmux_3_9_16153_16173 (
    .I(net_16153),
    .O(net_16173)
  );
  InMux inmux_3_9_16156_16179 (
    .I(net_16156),
    .O(net_16179)
  );
  InMux inmux_3_9_16158_16168 (
    .I(net_16158),
    .O(net_16168)
  );
  InMux inmux_3_9_16164_16174 (
    .I(net_16164),
    .O(net_16174)
  );
  InMux inmux_3_9_16170_16180 (
    .I(net_16170),
    .O(net_16180)
  );
  InMux inmux_3_9_16176_16186 (
    .I(net_16176),
    .O(net_16186)
  );
  InMux inmux_3_9_16182_16192 (
    .I(net_16182),
    .O(net_16192)
  );
  InMux inmux_3_9_16188_16198 (
    .I(net_16188),
    .O(net_16198)
  );
  InMux inmux_3_9_16194_16204 (
    .I(net_16194),
    .O(net_16204)
  );
  InMux inmux_4_10_20075_20116 (
    .I(net_20075),
    .O(net_20116)
  );
  InMux inmux_4_10_20101_20114 (
    .I(net_20101),
    .O(net_20114)
  );
  InMux inmux_4_10_20101_20121 (
    .I(net_20101),
    .O(net_20121)
  );
  InMux inmux_4_10_20101_20126 (
    .I(net_20101),
    .O(net_20126)
  );
  InMux inmux_4_10_20101_20133 (
    .I(net_20101),
    .O(net_20133)
  );
  InMux inmux_4_10_20101_20138 (
    .I(net_20101),
    .O(net_20138)
  );
  InMux inmux_4_10_20101_20145 (
    .I(net_20101),
    .O(net_20145)
  );
  InMux inmux_4_10_20101_20150 (
    .I(net_20101),
    .O(net_20150)
  );
  InMux inmux_4_10_20101_20155 (
    .I(net_20101),
    .O(net_20155)
  );
  InMux inmux_4_10_20111_20115 (
    .I(net_20111),
    .O(net_20115)
  );
  InMux inmux_4_10_20111_20120 (
    .I(net_20111),
    .O(net_20120)
  );
  InMux inmux_4_10_20111_20127 (
    .I(net_20111),
    .O(net_20127)
  );
  InMux inmux_4_10_20111_20132 (
    .I(net_20111),
    .O(net_20132)
  );
  InMux inmux_4_10_20111_20139 (
    .I(net_20111),
    .O(net_20139)
  );
  InMux inmux_4_10_20111_20144 (
    .I(net_20111),
    .O(net_20144)
  );
  InMux inmux_4_10_20111_20151 (
    .I(net_20111),
    .O(net_20151)
  );
  InMux inmux_4_10_20111_20156 (
    .I(net_20111),
    .O(net_20156)
  );
  InMux inmux_4_10_20112_20122 (
    .I(net_20112),
    .O(net_20122)
  );
  InMux inmux_4_10_20118_20128 (
    .I(net_20118),
    .O(net_20128)
  );
  InMux inmux_4_10_20124_20134 (
    .I(net_20124),
    .O(net_20134)
  );
  InMux inmux_4_10_20130_20140 (
    .I(net_20130),
    .O(net_20140)
  );
  InMux inmux_4_10_20136_20146 (
    .I(net_20136),
    .O(net_20146)
  );
  InMux inmux_4_10_20142_20152 (
    .I(net_20142),
    .O(net_20152)
  );
  InMux inmux_4_10_20148_20158 (
    .I(net_20148),
    .O(net_20158)
  );
  ClkMux inmux_4_10_5_20160 (
    .I(net_5),
    .O(net_20160)
  );
  SRMux inmux_4_10_9_20161 (
    .I(net_9),
    .O(net_20161)
  );
  InMux inmux_4_11_20204_20266 (
    .I(net_20204),
    .O(net_20266)
  );
  InMux inmux_4_11_20205_20281 (
    .I(net_20205),
    .O(net_20281)
  );
  InMux inmux_4_11_20207_20255 (
    .I(net_20207),
    .O(net_20255)
  );
  InMux inmux_4_11_20213_20251 (
    .I(net_20213),
    .O(net_20251)
  );
  InMux inmux_4_11_20215_20237 (
    .I(net_20215),
    .O(net_20237)
  );
  InMux inmux_4_11_20220_20242 (
    .I(net_20220),
    .O(net_20242)
  );
  InMux inmux_4_11_20228_20262 (
    .I(net_20228),
    .O(net_20262)
  );
  InMux inmux_4_11_20232_20274 (
    .I(net_20232),
    .O(net_20274)
  );
  ClkMux inmux_4_11_5_20283 (
    .I(net_5),
    .O(net_20283)
  );
  SRMux inmux_4_11_9_20284 (
    .I(net_9),
    .O(net_20284)
  );
  CEMux inmux_4_12_10_20405 (
    .I(net_10),
    .O(net_20405)
  );
  InMux inmux_4_12_20333_20391 (
    .I(net_20333),
    .O(net_20391)
  );
  InMux inmux_4_12_20337_20383 (
    .I(net_20337),
    .O(net_20383)
  );
  InMux inmux_4_12_20341_20380 (
    .I(net_20341),
    .O(net_20380)
  );
  InMux inmux_4_12_20344_20404 (
    .I(net_20344),
    .O(net_20404)
  );
  InMux inmux_4_12_20348_20371 (
    .I(net_20348),
    .O(net_20371)
  );
  InMux inmux_4_12_20350_20367 (
    .I(net_20350),
    .O(net_20367)
  );
  InMux inmux_4_12_20352_20362 (
    .I(net_20352),
    .O(net_20362)
  );
  ClkMux inmux_4_12_5_20406 (
    .I(net_5),
    .O(net_20406)
  );
  InMux inmux_4_13_20449_20501 (
    .I(net_20449),
    .O(net_20501)
  );
  InMux inmux_4_13_20450_20502 (
    .I(net_20450),
    .O(net_20502)
  );
  InMux inmux_4_13_20452_20495 (
    .I(net_20452),
    .O(net_20495)
  );
  InMux inmux_4_13_20453_20513 (
    .I(net_20453),
    .O(net_20513)
  );
  InMux inmux_4_13_20455_20484 (
    .I(net_20455),
    .O(net_20484)
  );
  InMux inmux_4_13_20459_20483 (
    .I(net_20459),
    .O(net_20483)
  );
  InMux inmux_4_13_20460_20520 (
    .I(net_20460),
    .O(net_20520)
  );
  InMux inmux_4_13_20466_20507 (
    .I(net_20466),
    .O(net_20507)
  );
  InMux inmux_4_13_20470_20514 (
    .I(net_20470),
    .O(net_20514)
  );
  InMux inmux_4_13_20471_20496 (
    .I(net_20471),
    .O(net_20496)
  );
  InMux inmux_4_13_20472_20519 (
    .I(net_20472),
    .O(net_20519)
  );
  InMux inmux_4_13_20476_20489 (
    .I(net_20476),
    .O(net_20489)
  );
  InMux inmux_4_13_20477_20490 (
    .I(net_20477),
    .O(net_20490)
  );
  InMux inmux_4_13_20478_20508 (
    .I(net_20478),
    .O(net_20508)
  );
  InMux inmux_4_13_20517_20527 (
    .I(net_20517),
    .O(net_20527)
  );
  InMux inmux_4_14_20584_20606 (
    .I(net_20584),
    .O(net_20606)
  );
  InMux inmux_4_14_20591_20611 (
    .I(net_20591),
    .O(net_20611)
  );
  InMux inmux_4_14_20593_20644 (
    .I(net_20593),
    .O(net_20644)
  );
  InMux inmux_4_14_20596_20647 (
    .I(net_20596),
    .O(net_20647)
  );
  InMux inmux_4_14_20598_20637 (
    .I(net_20598),
    .O(net_20637)
  );
  InMux inmux_4_14_20601_20629 (
    .I(net_20601),
    .O(net_20629)
  );
  InMux inmux_4_14_20602_20625 (
    .I(net_20602),
    .O(net_20625)
  );
  ClkMux inmux_4_14_5_20652 (
    .I(net_5),
    .O(net_20652)
  );
  SRMux inmux_4_14_9_20653 (
    .I(net_9),
    .O(net_20653)
  );
  InMux inmux_4_15_20695_20759 (
    .I(net_20695),
    .O(net_20759)
  );
  InMux inmux_4_15_20712_20746 (
    .I(net_20712),
    .O(net_20746)
  );
  InMux inmux_4_15_20713_20728 (
    .I(net_20713),
    .O(net_20728)
  );
  InMux inmux_4_15_20715_20752 (
    .I(net_20715),
    .O(net_20752)
  );
  InMux inmux_4_15_20717_20737 (
    .I(net_20717),
    .O(net_20737)
  );
  InMux inmux_4_15_20721_20770 (
    .I(net_20721),
    .O(net_20770)
  );
  InMux inmux_4_15_20725_20743 (
    .I(net_20725),
    .O(net_20743)
  );
  InMux inmux_4_15_20726_20766 (
    .I(net_20726),
    .O(net_20766)
  );
  ClkMux inmux_4_15_5_20775 (
    .I(net_5),
    .O(net_20775)
  );
  SRMux inmux_4_15_9_20776 (
    .I(net_9),
    .O(net_20776)
  );
  InMux inmux_4_16_20818_20858 (
    .I(net_20818),
    .O(net_20858)
  );
  InMux inmux_4_16_20825_20883 (
    .I(net_20825),
    .O(net_20883)
  );
  InMux inmux_4_16_20831_20877 (
    .I(net_20831),
    .O(net_20877)
  );
  InMux inmux_4_16_20834_20896 (
    .I(net_20834),
    .O(net_20896)
  );
  InMux inmux_4_16_20841_20852 (
    .I(net_20841),
    .O(net_20852)
  );
  InMux inmux_4_16_20846_20888 (
    .I(net_20846),
    .O(net_20888)
  );
  ClkMux inmux_4_16_5_20898 (
    .I(net_5),
    .O(net_20898)
  );
  SRMux inmux_4_16_9_20899 (
    .I(net_9),
    .O(net_20899)
  );
  InMux inmux_4_17_20942_21006 (
    .I(net_20942),
    .O(net_21006)
  );
  InMux inmux_4_17_20949_20980 (
    .I(net_20949),
    .O(net_20980)
  );
  InMux inmux_4_17_20952_21017 (
    .I(net_20952),
    .O(net_21017)
  );
  InMux inmux_4_17_20954_20993 (
    .I(net_20954),
    .O(net_20993)
  );
  InMux inmux_4_17_20955_21001 (
    .I(net_20955),
    .O(net_21001)
  );
  InMux inmux_4_17_20958_20977 (
    .I(net_20958),
    .O(net_20977)
  );
  InMux inmux_4_17_20967_21013 (
    .I(net_20967),
    .O(net_21013)
  );
  ClkMux inmux_4_17_5_21021 (
    .I(net_5),
    .O(net_21021)
  );
  SRMux inmux_4_17_9_21022 (
    .I(net_9),
    .O(net_21022)
  );
  InMux inmux_4_18_21070_21118 (
    .I(net_21070),
    .O(net_21118)
  );
  InMux inmux_4_18_21075_21116 (
    .I(net_21075),
    .O(net_21116)
  );
  InMux inmux_4_18_21078_21117 (
    .I(net_21078),
    .O(net_21117)
  );
  InMux inmux_4_18_21088_21115 (
    .I(net_21088),
    .O(net_21115)
  );
  CEMux inmux_4_18_21091_21143 (
    .I(net_21091),
    .O(net_21143)
  );
  ClkMux inmux_4_18_5_21144 (
    .I(net_5),
    .O(net_21144)
  );
  SRMux inmux_4_18_9_21145 (
    .I(net_9),
    .O(net_21145)
  );
  InMux inmux_4_19_21192_21264 (
    .I(net_21192),
    .O(net_21264)
  );
  InMux inmux_4_19_21196_21222 (
    .I(net_21196),
    .O(net_21222)
  );
  InMux inmux_4_19_21205_21258 (
    .I(net_21205),
    .O(net_21258)
  );
  ClkMux inmux_4_19_5_21267 (
    .I(net_5),
    .O(net_21267)
  );
  SRMux inmux_4_19_9_21268 (
    .I(net_9),
    .O(net_21268)
  );
  InMux inmux_4_1_18935_19011 (
    .I(net_18935),
    .O(net_19011)
  );
  InMux inmux_4_1_18936_19010 (
    .I(net_18936),
    .O(net_19010)
  );
  InMux inmux_4_1_18940_18969 (
    .I(net_18940),
    .O(net_18969)
  );
  InMux inmux_4_1_18942_18968 (
    .I(net_18942),
    .O(net_18968)
  );
  InMux inmux_4_1_18942_18985 (
    .I(net_18942),
    .O(net_18985)
  );
  InMux inmux_4_1_18942_18992 (
    .I(net_18942),
    .O(net_18992)
  );
  InMux inmux_4_1_18942_19002 (
    .I(net_18942),
    .O(net_19002)
  );
  InMux inmux_4_1_18942_19009 (
    .I(net_18942),
    .O(net_19009)
  );
  InMux inmux_4_1_18943_19005 (
    .I(net_18943),
    .O(net_19005)
  );
  InMux inmux_4_1_18944_19004 (
    .I(net_18944),
    .O(net_19004)
  );
  InMux inmux_4_1_18945_18996 (
    .I(net_18945),
    .O(net_18996)
  );
  InMux inmux_4_1_18946_18999 (
    .I(net_18946),
    .O(net_18999)
  );
  InMux inmux_4_1_18948_18966 (
    .I(net_18948),
    .O(net_18966)
  );
  InMux inmux_4_1_18949_18980 (
    .I(net_18949),
    .O(net_18980)
  );
  CEMux inmux_4_1_18951_19012 (
    .I(net_18951),
    .O(net_19012)
  );
  InMux inmux_4_1_18952_18967 (
    .I(net_18952),
    .O(net_18967)
  );
  InMux inmux_4_1_18952_18991 (
    .I(net_18952),
    .O(net_18991)
  );
  InMux inmux_4_1_18952_18998 (
    .I(net_18952),
    .O(net_18998)
  );
  InMux inmux_4_1_18952_19003 (
    .I(net_18952),
    .O(net_19003)
  );
  InMux inmux_4_1_18952_19008 (
    .I(net_18952),
    .O(net_19008)
  );
  InMux inmux_4_1_18954_18984 (
    .I(net_18954),
    .O(net_18984)
  );
  InMux inmux_4_1_18960_18978 (
    .I(net_18960),
    .O(net_18978)
  );
  InMux inmux_4_1_18960_18990 (
    .I(net_18960),
    .O(net_18990)
  );
  InMux inmux_4_1_18960_18997 (
    .I(net_18960),
    .O(net_18997)
  );
  InMux inmux_4_1_18963_18993 (
    .I(net_18963),
    .O(net_18993)
  );
  ClkMux inmux_4_1_5_19013 (
    .I(net_5),
    .O(net_19013)
  );
  SRMux inmux_4_1_9_19014 (
    .I(net_9),
    .O(net_19014)
  );
  InMux inmux_4_20_21315_21368 (
    .I(net_21315),
    .O(net_21368)
  );
  InMux inmux_4_20_21317_21375 (
    .I(net_21317),
    .O(net_21375)
  );
  ClkMux inmux_4_20_5_21390 (
    .I(net_5),
    .O(net_21390)
  );
  SRMux inmux_4_20_9_21391 (
    .I(net_9),
    .O(net_21391)
  );
  InMux inmux_4_22_21579_21626 (
    .I(net_21579),
    .O(net_21626)
  );
  ClkMux inmux_4_22_5_21636 (
    .I(net_5),
    .O(net_21636)
  );
  SRMux inmux_4_22_9_21637 (
    .I(net_9),
    .O(net_21637)
  );
  InMux inmux_4_2_19098_19155 (
    .I(net_19098),
    .O(net_19155)
  );
  InMux inmux_4_2_19100_19167 (
    .I(net_19100),
    .O(net_19167)
  );
  InMux inmux_4_2_19102_19131 (
    .I(net_19102),
    .O(net_19131)
  );
  InMux inmux_4_2_19103_19161 (
    .I(net_19103),
    .O(net_19161)
  );
  InMux inmux_4_2_19107_19172 (
    .I(net_19107),
    .O(net_19172)
  );
  InMux inmux_4_2_19108_19137 (
    .I(net_19108),
    .O(net_19137)
  );
  InMux inmux_4_2_19109_19136 (
    .I(net_19109),
    .O(net_19136)
  );
  InMux inmux_4_2_19110_19149 (
    .I(net_19110),
    .O(net_19149)
  );
  InMux inmux_4_2_19113_19166 (
    .I(net_19113),
    .O(net_19166)
  );
  InMux inmux_4_2_19114_19148 (
    .I(net_19114),
    .O(net_19148)
  );
  InMux inmux_4_2_19117_19142 (
    .I(net_19117),
    .O(net_19142)
  );
  InMux inmux_4_2_19118_19153 (
    .I(net_19118),
    .O(net_19153)
  );
  InMux inmux_4_2_19118_19165 (
    .I(net_19118),
    .O(net_19165)
  );
  InMux inmux_4_2_19119_19173 (
    .I(net_19119),
    .O(net_19173)
  );
  InMux inmux_4_2_19122_19130 (
    .I(net_19122),
    .O(net_19130)
  );
  InMux inmux_4_2_19123_19143 (
    .I(net_19123),
    .O(net_19143)
  );
  InMux inmux_4_2_19124_19154 (
    .I(net_19124),
    .O(net_19154)
  );
  InMux inmux_4_2_19126_19135 (
    .I(net_19126),
    .O(net_19135)
  );
  InMux inmux_4_2_19126_19159 (
    .I(net_19126),
    .O(net_19159)
  );
  InMux inmux_4_2_19127_19160 (
    .I(net_19127),
    .O(net_19160)
  );
  InMux inmux_4_2_19128_19138 (
    .I(net_19128),
    .O(net_19138)
  );
  InMux inmux_4_2_19134_19144 (
    .I(net_19134),
    .O(net_19144)
  );
  InMux inmux_4_2_19140_19150 (
    .I(net_19140),
    .O(net_19150)
  );
  InMux inmux_4_2_19146_19156 (
    .I(net_19146),
    .O(net_19156)
  );
  InMux inmux_4_2_19152_19162 (
    .I(net_19152),
    .O(net_19162)
  );
  InMux inmux_4_2_19158_19168 (
    .I(net_19158),
    .O(net_19168)
  );
  InMux inmux_4_2_19164_19174 (
    .I(net_19164),
    .O(net_19174)
  );
  InMux inmux_4_3_19214_19255 (
    .I(net_19214),
    .O(net_19255)
  );
  InMux inmux_4_3_19219_19259 (
    .I(net_19219),
    .O(net_19259)
  );
  InMux inmux_4_3_19221_19271 (
    .I(net_19221),
    .O(net_19271)
  );
  InMux inmux_4_3_19222_19265 (
    .I(net_19222),
    .O(net_19265)
  );
  InMux inmux_4_3_19223_19254 (
    .I(net_19223),
    .O(net_19254)
  );
  InMux inmux_4_3_19224_19260 (
    .I(net_19224),
    .O(net_19260)
  );
  InMux inmux_4_3_19225_19290 (
    .I(net_19225),
    .O(net_19290)
  );
  InMux inmux_4_3_19230_19252 (
    .I(net_19230),
    .O(net_19252)
  );
  InMux inmux_4_3_19230_19297 (
    .I(net_19230),
    .O(net_19297)
  );
  InMux inmux_4_3_19231_19296 (
    .I(net_19231),
    .O(net_19296)
  );
  InMux inmux_4_3_19232_19295 (
    .I(net_19232),
    .O(net_19295)
  );
  InMux inmux_4_3_19233_19272 (
    .I(net_19233),
    .O(net_19272)
  );
  InMux inmux_4_3_19233_19277 (
    .I(net_19233),
    .O(net_19277)
  );
  InMux inmux_4_3_19234_19285 (
    .I(net_19234),
    .O(net_19285)
  );
  InMux inmux_4_3_19236_19294 (
    .I(net_19236),
    .O(net_19294)
  );
  CEMux inmux_4_3_19237_19298 (
    .I(net_19237),
    .O(net_19298)
  );
  InMux inmux_4_3_19239_19266 (
    .I(net_19239),
    .O(net_19266)
  );
  InMux inmux_4_3_19240_19253 (
    .I(net_19240),
    .O(net_19253)
  );
  InMux inmux_4_3_19241_19276 (
    .I(net_19241),
    .O(net_19276)
  );
  InMux inmux_4_3_19242_19284 (
    .I(net_19242),
    .O(net_19284)
  );
  InMux inmux_4_3_19242_19289 (
    .I(net_19242),
    .O(net_19289)
  );
  InMux inmux_4_3_19245_19282 (
    .I(net_19245),
    .O(net_19282)
  );
  InMux inmux_4_3_19247_19291 (
    .I(net_19247),
    .O(net_19291)
  );
  InMux inmux_4_3_19250_19283 (
    .I(net_19250),
    .O(net_19283)
  );
  InMux inmux_4_3_19251_19261 (
    .I(net_19251),
    .O(net_19261)
  );
  InMux inmux_4_3_19257_19267 (
    .I(net_19257),
    .O(net_19267)
  );
  InMux inmux_4_3_19263_19273 (
    .I(net_19263),
    .O(net_19273)
  );
  InMux inmux_4_3_19269_19279 (
    .I(net_19269),
    .O(net_19279)
  );
  ClkMux inmux_4_3_5_19299 (
    .I(net_5),
    .O(net_19299)
  );
  SRMux inmux_4_3_9_19300 (
    .I(net_9),
    .O(net_19300)
  );
  InMux inmux_4_4_19346_19394 (
    .I(net_19346),
    .O(net_19394)
  );
  InMux inmux_4_4_19348_19384 (
    .I(net_19348),
    .O(net_19384)
  );
  InMux inmux_4_4_19350_19376 (
    .I(net_19350),
    .O(net_19376)
  );
  InMux inmux_4_4_19350_19395 (
    .I(net_19350),
    .O(net_19395)
  );
  InMux inmux_4_4_19352_19414 (
    .I(net_19352),
    .O(net_19414)
  );
  InMux inmux_4_4_19353_19399 (
    .I(net_19353),
    .O(net_19399)
  );
  InMux inmux_4_4_19354_19378 (
    .I(net_19354),
    .O(net_19378)
  );
  InMux inmux_4_4_19356_19402 (
    .I(net_19356),
    .O(net_19402)
  );
  InMux inmux_4_4_19356_19412 (
    .I(net_19356),
    .O(net_19412)
  );
  InMux inmux_4_4_19360_19408 (
    .I(net_19360),
    .O(net_19408)
  );
  InMux inmux_4_4_19361_19393 (
    .I(net_19361),
    .O(net_19393)
  );
  InMux inmux_4_4_19362_19413 (
    .I(net_19362),
    .O(net_19413)
  );
  InMux inmux_4_4_19365_19390 (
    .I(net_19365),
    .O(net_19390)
  );
  InMux inmux_4_4_19371_19401 (
    .I(net_19371),
    .O(net_19401)
  );
  InMux inmux_4_4_19373_19377 (
    .I(net_19373),
    .O(net_19377)
  );
  InMux inmux_4_4_19373_19396 (
    .I(net_19373),
    .O(net_19396)
  );
  InMux inmux_4_4_19373_19411 (
    .I(net_19373),
    .O(net_19411)
  );
  ClkMux inmux_4_4_5_19422 (
    .I(net_5),
    .O(net_19422)
  );
  SRMux inmux_4_4_9_19423 (
    .I(net_9),
    .O(net_19423)
  );
  InMux inmux_4_5_19470_19523 (
    .I(net_19470),
    .O(net_19523)
  );
  InMux inmux_4_5_19471_19519 (
    .I(net_19471),
    .O(net_19519)
  );
  InMux inmux_4_5_19473_19516 (
    .I(net_19473),
    .O(net_19516)
  );
  InMux inmux_4_5_19474_19500 (
    .I(net_19474),
    .O(net_19500)
  );
  InMux inmux_4_5_19478_19531 (
    .I(net_19478),
    .O(net_19531)
  );
  InMux inmux_4_5_19479_19525 (
    .I(net_19479),
    .O(net_19525)
  );
  InMux inmux_4_5_19479_19530 (
    .I(net_19479),
    .O(net_19530)
  );
  InMux inmux_4_5_19481_19524 (
    .I(net_19481),
    .O(net_19524)
  );
  InMux inmux_4_5_19481_19529 (
    .I(net_19481),
    .O(net_19529)
  );
  InMux inmux_4_5_19483_19536 (
    .I(net_19483),
    .O(net_19536)
  );
  InMux inmux_4_5_19485_19534 (
    .I(net_19485),
    .O(net_19534)
  );
  InMux inmux_4_5_19488_19513 (
    .I(net_19488),
    .O(net_19513)
  );
  InMux inmux_4_5_19492_19498 (
    .I(net_19492),
    .O(net_19498)
  );
  InMux inmux_4_5_19493_19535 (
    .I(net_19493),
    .O(net_19535)
  );
  InMux inmux_4_5_19494_19541 (
    .I(net_19494),
    .O(net_19541)
  );
  InMux inmux_4_5_19495_19537 (
    .I(net_19495),
    .O(net_19537)
  );
  InMux inmux_4_5_19496_19505 (
    .I(net_19496),
    .O(net_19505)
  );
  ClkMux inmux_4_5_5_19545 (
    .I(net_5),
    .O(net_19545)
  );
  SRMux inmux_4_5_9_19546 (
    .I(net_9),
    .O(net_19546)
  );
  InMux inmux_4_6_19588_19647 (
    .I(net_19588),
    .O(net_19647)
  );
  InMux inmux_4_6_19590_19659 (
    .I(net_19590),
    .O(net_19659)
  );
  InMux inmux_4_6_19591_19627 (
    .I(net_19591),
    .O(net_19627)
  );
  InMux inmux_4_6_19592_19623 (
    .I(net_19592),
    .O(net_19623)
  );
  InMux inmux_4_6_19595_19648 (
    .I(net_19595),
    .O(net_19648)
  );
  InMux inmux_4_6_19596_19646 (
    .I(net_19596),
    .O(net_19646)
  );
  InMux inmux_4_6_19599_19633 (
    .I(net_19599),
    .O(net_19633)
  );
  InMux inmux_4_6_19602_19651 (
    .I(net_19602),
    .O(net_19651)
  );
  InMux inmux_4_6_19603_19642 (
    .I(net_19603),
    .O(net_19642)
  );
  InMux inmux_4_6_19604_19664 (
    .I(net_19604),
    .O(net_19664)
  );
  InMux inmux_4_6_19612_19629 (
    .I(net_19612),
    .O(net_19629)
  );
  InMux inmux_4_6_19612_19636 (
    .I(net_19612),
    .O(net_19636)
  );
  InMux inmux_4_6_19612_19641 (
    .I(net_19612),
    .O(net_19641)
  );
  InMux inmux_4_6_19612_19653 (
    .I(net_19612),
    .O(net_19653)
  );
  InMux inmux_4_6_19612_19660 (
    .I(net_19612),
    .O(net_19660)
  );
  InMux inmux_4_6_19615_19645 (
    .I(net_19615),
    .O(net_19645)
  );
  ClkMux inmux_4_6_5_19668 (
    .I(net_5),
    .O(net_19668)
  );
  CEMux inmux_4_6_8_19667 (
    .I(net_8),
    .O(net_19667)
  );
  InMux inmux_4_7_19712_19769 (
    .I(net_19712),
    .O(net_19769)
  );
  InMux inmux_4_7_19715_19765 (
    .I(net_19715),
    .O(net_19765)
  );
  InMux inmux_4_7_19718_19757 (
    .I(net_19718),
    .O(net_19757)
  );
  InMux inmux_4_7_19720_19763 (
    .I(net_19720),
    .O(net_19763)
  );
  InMux inmux_4_7_19721_19762 (
    .I(net_19721),
    .O(net_19762)
  );
  InMux inmux_4_7_19721_19771 (
    .I(net_19721),
    .O(net_19771)
  );
  InMux inmux_4_7_19724_19780 (
    .I(net_19724),
    .O(net_19780)
  );
  InMux inmux_4_7_19725_19745 (
    .I(net_19725),
    .O(net_19745)
  );
  InMux inmux_4_7_19726_19758 (
    .I(net_19726),
    .O(net_19758)
  );
  InMux inmux_4_7_19729_19768 (
    .I(net_19729),
    .O(net_19768)
  );
  InMux inmux_4_7_19731_19753 (
    .I(net_19731),
    .O(net_19753)
  );
  InMux inmux_4_7_19732_19788 (
    .I(net_19732),
    .O(net_19788)
  );
  InMux inmux_4_7_19734_19759 (
    .I(net_19734),
    .O(net_19759)
  );
  InMux inmux_4_7_19735_19764 (
    .I(net_19735),
    .O(net_19764)
  );
  InMux inmux_4_7_19736_19746 (
    .I(net_19736),
    .O(net_19746)
  );
  InMux inmux_4_7_19736_19756 (
    .I(net_19736),
    .O(net_19756)
  );
  InMux inmux_4_7_19737_19747 (
    .I(net_19737),
    .O(net_19747)
  );
  InMux inmux_4_7_19738_19770 (
    .I(net_19738),
    .O(net_19770)
  );
  InMux inmux_4_7_19740_19744 (
    .I(net_19740),
    .O(net_19744)
  );
  InMux inmux_4_7_19742_19775 (
    .I(net_19742),
    .O(net_19775)
  );
  ClkMux inmux_4_7_5_19791 (
    .I(net_5),
    .O(net_19791)
  );
  CEMux inmux_4_7_8_19790 (
    .I(net_8),
    .O(net_19790)
  );
  InMux inmux_4_8_19838_19869 (
    .I(net_19838),
    .O(net_19869)
  );
  InMux inmux_4_8_19848_19868 (
    .I(net_19848),
    .O(net_19868)
  );
  InMux inmux_4_8_19848_19875 (
    .I(net_19848),
    .O(net_19875)
  );
  InMux inmux_4_8_19848_19880 (
    .I(net_19848),
    .O(net_19880)
  );
  InMux inmux_4_8_19848_19887 (
    .I(net_19848),
    .O(net_19887)
  );
  InMux inmux_4_8_19848_19892 (
    .I(net_19848),
    .O(net_19892)
  );
  InMux inmux_4_8_19848_19899 (
    .I(net_19848),
    .O(net_19899)
  );
  InMux inmux_4_8_19848_19904 (
    .I(net_19848),
    .O(net_19904)
  );
  InMux inmux_4_8_19848_19911 (
    .I(net_19848),
    .O(net_19911)
  );
  InMux inmux_4_8_19852_19881 (
    .I(net_19852),
    .O(net_19881)
  );
  InMux inmux_4_8_19854_19893 (
    .I(net_19854),
    .O(net_19893)
  );
  InMux inmux_4_8_19856_19905 (
    .I(net_19856),
    .O(net_19905)
  );
  InMux inmux_4_8_19859_19874 (
    .I(net_19859),
    .O(net_19874)
  );
  InMux inmux_4_8_19861_19886 (
    .I(net_19861),
    .O(net_19886)
  );
  InMux inmux_4_8_19863_19898 (
    .I(net_19863),
    .O(net_19898)
  );
  InMux inmux_4_8_19865_19910 (
    .I(net_19865),
    .O(net_19910)
  );
  InMux inmux_4_8_19902_19912 (
    .I(net_19902),
    .O(net_19912)
  );
  ClkMux inmux_4_8_5_19914 (
    .I(net_5),
    .O(net_19914)
  );
  SRMux inmux_4_8_9_19915 (
    .I(net_9),
    .O(net_19915)
  );
  InMux inmux_4_9_19952_19993 (
    .I(net_19952),
    .O(net_19993)
  );
  InMux inmux_4_9_19960_19991 (
    .I(net_19960),
    .O(net_19991)
  );
  InMux inmux_4_9_19960_19998 (
    .I(net_19960),
    .O(net_19998)
  );
  InMux inmux_4_9_19960_20003 (
    .I(net_19960),
    .O(net_20003)
  );
  InMux inmux_4_9_19960_20010 (
    .I(net_19960),
    .O(net_20010)
  );
  InMux inmux_4_9_19960_20015 (
    .I(net_19960),
    .O(net_20015)
  );
  InMux inmux_4_9_19960_20022 (
    .I(net_19960),
    .O(net_20022)
  );
  InMux inmux_4_9_19960_20027 (
    .I(net_19960),
    .O(net_20027)
  );
  InMux inmux_4_9_19960_20034 (
    .I(net_19960),
    .O(net_20034)
  );
  InMux inmux_4_9_19972_19992 (
    .I(net_19972),
    .O(net_19992)
  );
  InMux inmux_4_9_19972_19997 (
    .I(net_19972),
    .O(net_19997)
  );
  InMux inmux_4_9_19972_20004 (
    .I(net_19972),
    .O(net_20004)
  );
  InMux inmux_4_9_19972_20009 (
    .I(net_19972),
    .O(net_20009)
  );
  InMux inmux_4_9_19972_20016 (
    .I(net_19972),
    .O(net_20016)
  );
  InMux inmux_4_9_19972_20021 (
    .I(net_19972),
    .O(net_20021)
  );
  InMux inmux_4_9_19972_20028 (
    .I(net_19972),
    .O(net_20028)
  );
  InMux inmux_4_9_19972_20033 (
    .I(net_19972),
    .O(net_20033)
  );
  InMux inmux_4_9_19989_19999 (
    .I(net_19989),
    .O(net_19999)
  );
  InMux inmux_4_9_19995_20005 (
    .I(net_19995),
    .O(net_20005)
  );
  InMux inmux_4_9_20001_20011 (
    .I(net_20001),
    .O(net_20011)
  );
  InMux inmux_4_9_20007_20017 (
    .I(net_20007),
    .O(net_20017)
  );
  InMux inmux_4_9_20013_20023 (
    .I(net_20013),
    .O(net_20023)
  );
  InMux inmux_4_9_20019_20029 (
    .I(net_20019),
    .O(net_20029)
  );
  InMux inmux_4_9_20025_20035 (
    .I(net_20025),
    .O(net_20035)
  );
  ClkMux inmux_4_9_5_20037 (
    .I(net_5),
    .O(net_20037)
  );
  SRMux inmux_4_9_9_20038 (
    .I(net_9),
    .O(net_20038)
  );
  IoInMux inmux_5_0_22721_22697 (
    .I(net_22721),
    .O(net_22697)
  );
  CEMux inmux_5_10_12_23990 (
    .I(net_12),
    .O(net_23990)
  );
  InMux inmux_5_10_23914_23947 (
    .I(net_23914),
    .O(net_23947)
  );
  InMux inmux_5_10_23916_23986 (
    .I(net_23916),
    .O(net_23986)
  );
  InMux inmux_5_10_23918_23981 (
    .I(net_23918),
    .O(net_23981)
  );
  InMux inmux_5_10_23920_23956 (
    .I(net_23920),
    .O(net_23956)
  );
  InMux inmux_5_10_23929_23953 (
    .I(net_23929),
    .O(net_23953)
  );
  InMux inmux_5_10_23933_23968 (
    .I(net_23933),
    .O(net_23968)
  );
  InMux inmux_5_10_23937_23974 (
    .I(net_23937),
    .O(net_23974)
  );
  InMux inmux_5_10_23939_23964 (
    .I(net_23939),
    .O(net_23964)
  );
  ClkMux inmux_5_10_5_23991 (
    .I(net_5),
    .O(net_23991)
  );
  InMux inmux_5_11_24042_24087 (
    .I(net_24042),
    .O(net_24087)
  );
  InMux inmux_5_11_24049_24074 (
    .I(net_24049),
    .O(net_24074)
  );
  InMux inmux_5_11_24050_24081 (
    .I(net_24050),
    .O(net_24081)
  );
  InMux inmux_5_11_24052_24067 (
    .I(net_24052),
    .O(net_24067)
  );
  InMux inmux_5_11_24054_24098 (
    .I(net_24054),
    .O(net_24098)
  );
  InMux inmux_5_11_24058_24109 (
    .I(net_24058),
    .O(net_24109)
  );
  InMux inmux_5_11_24060_24092 (
    .I(net_24060),
    .O(net_24092)
  );
  InMux inmux_5_11_24062_24104 (
    .I(net_24062),
    .O(net_24104)
  );
  ClkMux inmux_5_11_5_24114 (
    .I(net_5),
    .O(net_24114)
  );
  SRMux inmux_5_11_9_24115 (
    .I(net_9),
    .O(net_24115)
  );
  InMux inmux_5_12_24161_24199 (
    .I(net_24161),
    .O(net_24199)
  );
  InMux inmux_5_12_24164_24193 (
    .I(net_24164),
    .O(net_24193)
  );
  InMux inmux_5_12_24170_24235 (
    .I(net_24170),
    .O(net_24235)
  );
  InMux inmux_5_12_24173_24202 (
    .I(net_24173),
    .O(net_24202)
  );
  InMux inmux_5_12_24175_24216 (
    .I(net_24175),
    .O(net_24216)
  );
  InMux inmux_5_12_24177_24221 (
    .I(net_24177),
    .O(net_24221)
  );
  InMux inmux_5_12_24182_24226 (
    .I(net_24182),
    .O(net_24226)
  );
  InMux inmux_5_12_24184_24211 (
    .I(net_24184),
    .O(net_24211)
  );
  ClkMux inmux_5_12_5_24237 (
    .I(net_5),
    .O(net_24237)
  );
  SRMux inmux_5_12_9_24238 (
    .I(net_9),
    .O(net_24238)
  );
  InMux inmux_5_13_24283_24328 (
    .I(net_24283),
    .O(net_24328)
  );
  InMux inmux_5_13_24286_24320 (
    .I(net_24286),
    .O(net_24320)
  );
  InMux inmux_5_13_24293_24313 (
    .I(net_24293),
    .O(net_24313)
  );
  InMux inmux_5_13_24296_24344 (
    .I(net_24296),
    .O(net_24344)
  );
  InMux inmux_5_13_24298_24358 (
    .I(net_24298),
    .O(net_24358)
  );
  InMux inmux_5_13_24300_24337 (
    .I(net_24300),
    .O(net_24337)
  );
  InMux inmux_5_13_24306_24333 (
    .I(net_24306),
    .O(net_24333)
  );
  InMux inmux_5_13_24310_24350 (
    .I(net_24310),
    .O(net_24350)
  );
  ClkMux inmux_5_13_5_24360 (
    .I(net_5),
    .O(net_24360)
  );
  SRMux inmux_5_13_9_24361 (
    .I(net_9),
    .O(net_24361)
  );
  InMux inmux_5_14_24416_24443 (
    .I(net_24416),
    .O(net_24443)
  );
  InMux inmux_5_14_24421_24469 (
    .I(net_24421),
    .O(net_24469)
  );
  InMux inmux_5_14_24423_24438 (
    .I(net_24423),
    .O(net_24438)
  );
  InMux inmux_5_14_24428_24462 (
    .I(net_24428),
    .O(net_24462)
  );
  InMux inmux_5_14_24431_24451 (
    .I(net_24431),
    .O(net_24451)
  );
  InMux inmux_5_14_24432_24479 (
    .I(net_24432),
    .O(net_24479)
  );
  ClkMux inmux_5_14_5_24483 (
    .I(net_5),
    .O(net_24483)
  );
  SRMux inmux_5_14_9_24484 (
    .I(net_9),
    .O(net_24484)
  );
  InMux inmux_5_15_24533_24601 (
    .I(net_24533),
    .O(net_24601)
  );
  InMux inmux_5_15_24535_24566 (
    .I(net_24535),
    .O(net_24566)
  );
  InMux inmux_5_15_24538_24598 (
    .I(net_24538),
    .O(net_24598)
  );
  InMux inmux_5_15_24548_24571 (
    .I(net_24548),
    .O(net_24571)
  );
  InMux inmux_5_15_24551_24578 (
    .I(net_24551),
    .O(net_24578)
  );
  InMux inmux_5_15_24553_24583 (
    .I(net_24553),
    .O(net_24583)
  );
  InMux inmux_5_15_24557_24590 (
    .I(net_24557),
    .O(net_24590)
  );
  ClkMux inmux_5_15_5_24606 (
    .I(net_5),
    .O(net_24606)
  );
  SRMux inmux_5_15_9_24607 (
    .I(net_9),
    .O(net_24607)
  );
  InMux inmux_5_16_24649_24720 (
    .I(net_24649),
    .O(net_24720)
  );
  CEMux inmux_5_16_24651_24728 (
    .I(net_24651),
    .O(net_24728)
  );
  InMux inmux_5_16_24653_24715 (
    .I(net_24653),
    .O(net_24715)
  );
  InMux inmux_5_16_24654_24712 (
    .I(net_24654),
    .O(net_24712)
  );
  InMux inmux_5_16_24656_24726 (
    .I(net_24656),
    .O(net_24726)
  );
  InMux inmux_5_16_24657_24695 (
    .I(net_24657),
    .O(net_24695)
  );
  InMux inmux_5_16_24657_24714 (
    .I(net_24657),
    .O(net_24714)
  );
  InMux inmux_5_16_24657_24724 (
    .I(net_24657),
    .O(net_24724)
  );
  InMux inmux_5_16_24658_24718 (
    .I(net_24658),
    .O(net_24718)
  );
  InMux inmux_5_16_24659_24697 (
    .I(net_24659),
    .O(net_24697)
  );
  InMux inmux_5_16_24660_24727 (
    .I(net_24660),
    .O(net_24727)
  );
  InMux inmux_5_16_24661_24719 (
    .I(net_24661),
    .O(net_24719)
  );
  InMux inmux_5_16_24662_24725 (
    .I(net_24662),
    .O(net_24725)
  );
  InMux inmux_5_16_24665_24694 (
    .I(net_24665),
    .O(net_24694)
  );
  InMux inmux_5_16_24675_24721 (
    .I(net_24675),
    .O(net_24721)
  );
  InMux inmux_5_16_24676_24696 (
    .I(net_24676),
    .O(net_24696)
  );
  InMux inmux_5_16_24680_24713 (
    .I(net_24680),
    .O(net_24713)
  );
  ClkMux inmux_5_16_5_24729 (
    .I(net_5),
    .O(net_24729)
  );
  SRMux inmux_5_16_9_24730 (
    .I(net_9),
    .O(net_24730)
  );
  InMux inmux_5_17_24772_24812 (
    .I(net_24772),
    .O(net_24812)
  );
  InMux inmux_5_17_24773_24813 (
    .I(net_24773),
    .O(net_24813)
  );
  InMux inmux_5_17_24780_24811 (
    .I(net_24780),
    .O(net_24811)
  );
  CEMux inmux_5_17_24783_24851 (
    .I(net_24783),
    .O(net_24851)
  );
  InMux inmux_5_17_24792_24814 (
    .I(net_24792),
    .O(net_24814)
  );
  ClkMux inmux_5_17_5_24852 (
    .I(net_5),
    .O(net_24852)
  );
  SRMux inmux_5_17_9_24853 (
    .I(net_9),
    .O(net_24853)
  );
  CEMux inmux_5_18_10_24974 (
    .I(net_10),
    .O(net_24974)
  );
  InMux inmux_5_18_24895_24952 (
    .I(net_24895),
    .O(net_24952)
  );
  InMux inmux_5_18_24899_24937 (
    .I(net_24899),
    .O(net_24937)
  );
  InMux inmux_5_18_24925_24948 (
    .I(net_24925),
    .O(net_24948)
  );
  ClkMux inmux_5_18_5_24975 (
    .I(net_5),
    .O(net_24975)
  );
  InMux inmux_5_19_25024_25053 (
    .I(net_25024),
    .O(net_25053)
  );
  InMux inmux_5_19_25038_25077 (
    .I(net_25038),
    .O(net_25077)
  );
  ClkMux inmux_5_19_5_25098 (
    .I(net_5),
    .O(net_25098)
  );
  SRMux inmux_5_19_9_25099 (
    .I(net_9),
    .O(net_25099)
  );
  InMux inmux_5_1_22785_22817 (
    .I(net_22785),
    .O(net_22817)
  );
  InMux inmux_5_1_22785_22841 (
    .I(net_22785),
    .O(net_22841)
  );
  InMux inmux_5_1_22790_22815 (
    .I(net_22790),
    .O(net_22815)
  );
  InMux inmux_5_1_22791_22818 (
    .I(net_22791),
    .O(net_22818)
  );
  ClkMux inmux_5_1_5_22844 (
    .I(net_5),
    .O(net_22844)
  );
  SRMux inmux_5_1_9_22845 (
    .I(net_9),
    .O(net_22845)
  );
  InMux inmux_5_2_22944_22968 (
    .I(net_22944),
    .O(net_22968)
  );
  InMux inmux_5_2_22955_22990 (
    .I(net_22955),
    .O(net_22990)
  );
  ClkMux inmux_5_2_5_23007 (
    .I(net_5),
    .O(net_23007)
  );
  CEMux inmux_5_2_8_23006 (
    .I(net_8),
    .O(net_23006)
  );
  InMux inmux_5_3_23055_23125 (
    .I(net_23055),
    .O(net_23125)
  );
  InMux inmux_5_3_23056_23095 (
    .I(net_23056),
    .O(net_23095)
  );
  InMux inmux_5_3_23061_23126 (
    .I(net_23061),
    .O(net_23126)
  );
  InMux inmux_5_3_23063_23128 (
    .I(net_23063),
    .O(net_23128)
  );
  InMux inmux_5_3_23069_23113 (
    .I(net_23069),
    .O(net_23113)
  );
  InMux inmux_5_3_23071_23127 (
    .I(net_23071),
    .O(net_23127)
  );
  CEMux inmux_5_3_23077_23129 (
    .I(net_23077),
    .O(net_23129)
  );
  InMux inmux_5_3_23078_23108 (
    .I(net_23078),
    .O(net_23108)
  );
  ClkMux inmux_5_3_5_23130 (
    .I(net_5),
    .O(net_23130)
  );
  InMux inmux_5_4_23177_23220 (
    .I(net_23177),
    .O(net_23220)
  );
  InMux inmux_5_4_23179_23206 (
    .I(net_23179),
    .O(net_23206)
  );
  InMux inmux_5_4_23186_23232 (
    .I(net_23186),
    .O(net_23232)
  );
  InMux inmux_5_4_23188_23215 (
    .I(net_23188),
    .O(net_23215)
  );
  InMux inmux_5_4_23189_23237 (
    .I(net_23189),
    .O(net_23237)
  );
  InMux inmux_5_4_23190_23243 (
    .I(net_23190),
    .O(net_23243)
  );
  InMux inmux_5_4_23197_23224 (
    .I(net_23197),
    .O(net_23224)
  );
  InMux inmux_5_4_23198_23225 (
    .I(net_23198),
    .O(net_23225)
  );
  InMux inmux_5_4_23204_23251 (
    .I(net_23204),
    .O(net_23251)
  );
  ClkMux inmux_5_4_5_23253 (
    .I(net_5),
    .O(net_23253)
  );
  SRMux inmux_5_4_9_23254 (
    .I(net_9),
    .O(net_23254)
  );
  InMux inmux_5_5_23299_23330 (
    .I(net_23299),
    .O(net_23330)
  );
  InMux inmux_5_5_23301_23361 (
    .I(net_23301),
    .O(net_23361)
  );
  InMux inmux_5_5_23305_23336 (
    .I(net_23305),
    .O(net_23336)
  );
  InMux inmux_5_5_23306_23342 (
    .I(net_23306),
    .O(net_23342)
  );
  InMux inmux_5_5_23307_23348 (
    .I(net_23307),
    .O(net_23348)
  );
  InMux inmux_5_5_23308_23354 (
    .I(net_23308),
    .O(net_23354)
  );
  InMux inmux_5_5_23310_23366 (
    .I(net_23310),
    .O(net_23366)
  );
  InMux inmux_5_5_23327_23331 (
    .I(net_23327),
    .O(net_23331)
  );
  InMux inmux_5_5_23328_23338 (
    .I(net_23328),
    .O(net_23338)
  );
  InMux inmux_5_5_23334_23344 (
    .I(net_23334),
    .O(net_23344)
  );
  InMux inmux_5_5_23340_23350 (
    .I(net_23340),
    .O(net_23350)
  );
  InMux inmux_5_5_23346_23356 (
    .I(net_23346),
    .O(net_23356)
  );
  InMux inmux_5_5_23352_23362 (
    .I(net_23352),
    .O(net_23362)
  );
  InMux inmux_5_5_23358_23368 (
    .I(net_23358),
    .O(net_23368)
  );
  InMux inmux_5_5_23364_23374 (
    .I(net_23364),
    .O(net_23374)
  );
  ClkMux inmux_5_5_5_23376 (
    .I(net_5),
    .O(net_23376)
  );
  SRMux inmux_5_5_9_23377 (
    .I(net_9),
    .O(net_23377)
  );
  CEMux inmux_5_6_12_23498 (
    .I(net_12),
    .O(net_23498)
  );
  InMux inmux_5_6_23419_23478 (
    .I(net_23419),
    .O(net_23478)
  );
  InMux inmux_5_6_23421_23466 (
    .I(net_23421),
    .O(net_23466)
  );
  InMux inmux_5_6_23422_23484 (
    .I(net_23422),
    .O(net_23484)
  );
  InMux inmux_5_6_23423_23483 (
    .I(net_23423),
    .O(net_23483)
  );
  InMux inmux_5_6_23424_23465 (
    .I(net_23424),
    .O(net_23465)
  );
  InMux inmux_5_6_23425_23471 (
    .I(net_23425),
    .O(net_23471)
  );
  InMux inmux_5_6_23426_23477 (
    .I(net_23426),
    .O(net_23477)
  );
  InMux inmux_5_6_23427_23472 (
    .I(net_23427),
    .O(net_23472)
  );
  InMux inmux_5_6_23436_23496 (
    .I(net_23436),
    .O(net_23496)
  );
  InMux inmux_5_6_23443_23453 (
    .I(net_23443),
    .O(net_23453)
  );
  InMux inmux_5_6_23445_23460 (
    .I(net_23445),
    .O(net_23460)
  );
  InMux inmux_5_6_23446_23459 (
    .I(net_23446),
    .O(net_23459)
  );
  InMux inmux_5_6_23448_23454 (
    .I(net_23448),
    .O(net_23454)
  );
  InMux inmux_5_6_23451_23461 (
    .I(net_23451),
    .O(net_23461)
  );
  InMux inmux_5_6_23457_23467 (
    .I(net_23457),
    .O(net_23467)
  );
  InMux inmux_5_6_23463_23473 (
    .I(net_23463),
    .O(net_23473)
  );
  InMux inmux_5_6_23469_23479 (
    .I(net_23469),
    .O(net_23479)
  );
  InMux inmux_5_6_23475_23485 (
    .I(net_23475),
    .O(net_23485)
  );
  InMux inmux_5_6_23481_23491 (
    .I(net_23481),
    .O(net_23491)
  );
  ClkMux inmux_5_6_5_23499 (
    .I(net_5),
    .O(net_23499)
  );
  CEMux inmux_5_7_10_23621 (
    .I(net_10),
    .O(net_23621)
  );
  InMux inmux_5_7_23547_23583 (
    .I(net_23547),
    .O(net_23583)
  );
  InMux inmux_5_7_23547_23595 (
    .I(net_23547),
    .O(net_23595)
  );
  InMux inmux_5_7_23547_23605 (
    .I(net_23547),
    .O(net_23605)
  );
  InMux inmux_5_7_23548_23606 (
    .I(net_23548),
    .O(net_23606)
  );
  InMux inmux_5_7_23551_23608 (
    .I(net_23551),
    .O(net_23608)
  );
  InMux inmux_5_7_23553_23594 (
    .I(net_23553),
    .O(net_23594)
  );
  InMux inmux_5_7_23554_23607 (
    .I(net_23554),
    .O(net_23607)
  );
  InMux inmux_5_7_23555_23582 (
    .I(net_23555),
    .O(net_23582)
  );
  InMux inmux_5_7_23556_23581 (
    .I(net_23556),
    .O(net_23581)
  );
  InMux inmux_5_7_23556_23593 (
    .I(net_23556),
    .O(net_23593)
  );
  InMux inmux_5_7_23567_23589 (
    .I(net_23567),
    .O(net_23589)
  );
  InMux inmux_5_7_23571_23584 (
    .I(net_23571),
    .O(net_23584)
  );
  ClkMux inmux_5_7_5_23622 (
    .I(net_5),
    .O(net_23622)
  );
  InMux inmux_5_8_23668_23704 (
    .I(net_23668),
    .O(net_23704)
  );
  InMux inmux_5_8_23670_23728 (
    .I(net_23670),
    .O(net_23728)
  );
  InMux inmux_5_8_23671_23700 (
    .I(net_23671),
    .O(net_23700)
  );
  InMux inmux_5_8_23672_23706 (
    .I(net_23672),
    .O(net_23706)
  );
  InMux inmux_5_8_23674_23736 (
    .I(net_23674),
    .O(net_23736)
  );
  InMux inmux_5_8_23676_23719 (
    .I(net_23676),
    .O(net_23719)
  );
  InMux inmux_5_8_23678_23722 (
    .I(net_23678),
    .O(net_23722)
  );
  InMux inmux_5_8_23682_23711 (
    .I(net_23682),
    .O(net_23711)
  );
  InMux inmux_5_8_23684_23716 (
    .I(net_23684),
    .O(net_23716)
  );
  InMux inmux_5_8_23687_23741 (
    .I(net_23687),
    .O(net_23741)
  );
  ClkMux inmux_5_8_5_23745 (
    .I(net_5),
    .O(net_23745)
  );
  SRMux inmux_5_8_9_23746 (
    .I(net_9),
    .O(net_23746)
  );
  InMux inmux_5_9_23804_23842 (
    .I(net_23804),
    .O(net_23842)
  );
  InMux inmux_5_9_23805_23851 (
    .I(net_23805),
    .O(net_23851)
  );
  InMux inmux_5_9_23806_23828 (
    .I(net_23806),
    .O(net_23828)
  );
  InMux inmux_5_9_23807_23834 (
    .I(net_23807),
    .O(net_23834)
  );
  InMux inmux_5_9_23811_23848 (
    .I(net_23811),
    .O(net_23848)
  );
  InMux inmux_5_9_23812_23822 (
    .I(net_23812),
    .O(net_23822)
  );
  InMux inmux_5_9_23814_23860 (
    .I(net_23814),
    .O(net_23860)
  );
  InMux inmux_5_9_23817_23866 (
    .I(net_23817),
    .O(net_23866)
  );
  ClkMux inmux_5_9_5_23868 (
    .I(net_5),
    .O(net_23868)
  );
  SRMux inmux_5_9_9_23869 (
    .I(net_9),
    .O(net_23869)
  );
  CEMux inmux_6_10_27569_27611 (
    .I(net_27569),
    .O(net_27611)
  );
  ClkMux inmux_6_10_5_27610 (
    .I(net_5),
    .O(net_27610)
  );
  CEMux inmux_6_11_27655_27713 (
    .I(net_27655),
    .O(net_27713)
  );
  SRMux inmux_6_11_27657_27714 (
    .I(net_27657),
    .O(net_27714)
  );
  InMux inmux_6_11_27659_27702 (
    .I(net_27659),
    .O(net_27702)
  );
  InMux inmux_6_11_27665_27701 (
    .I(net_27665),
    .O(net_27701)
  );
  ClkMux inmux_6_11_5_27712 (
    .I(net_5),
    .O(net_27712)
  );
  CEMux inmux_6_12_27766_27815 (
    .I(net_27766),
    .O(net_27815)
  );
  ClkMux inmux_6_12_5_27814 (
    .I(net_5),
    .O(net_27814)
  );
  InMux inmux_6_3_26839_26877 (
    .I(net_26839),
    .O(net_26877)
  );
  InMux inmux_6_3_26839_26883 (
    .I(net_26839),
    .O(net_26883)
  );
  InMux inmux_6_3_26841_26891 (
    .I(net_26841),
    .O(net_26891)
  );
  InMux inmux_6_3_26843_26905 (
    .I(net_26843),
    .O(net_26905)
  );
  InMux inmux_6_3_26844_26885 (
    .I(net_26844),
    .O(net_26885)
  );
  InMux inmux_6_3_26847_26878 (
    .I(net_26847),
    .O(net_26878)
  );
  InMux inmux_6_3_26847_26884 (
    .I(net_26847),
    .O(net_26884)
  );
  InMux inmux_6_3_26849_26890 (
    .I(net_26849),
    .O(net_26890)
  );
  InMux inmux_6_3_26850_26886 (
    .I(net_26850),
    .O(net_26886)
  );
  InMux inmux_6_3_26853_26889 (
    .I(net_26853),
    .O(net_26889)
  );
  CEMux inmux_6_3_26855_26897 (
    .I(net_26855),
    .O(net_26897)
  );
  InMux inmux_6_3_26856_26906 (
    .I(net_26856),
    .O(net_26906)
  );
  InMux inmux_6_3_26860_26888 (
    .I(net_26860),
    .O(net_26888)
  );
  InMux inmux_6_3_26861_26880 (
    .I(net_26861),
    .O(net_26880)
  );
  InMux inmux_6_3_26861_26882 (
    .I(net_26861),
    .O(net_26882)
  );
  InMux inmux_6_3_26862_26899 (
    .I(net_26862),
    .O(net_26899)
  );
  InMux inmux_6_3_26866_26879 (
    .I(net_26866),
    .O(net_26879)
  );
  InMux inmux_6_3_26866_26881 (
    .I(net_26866),
    .O(net_26881)
  );
  SRMux inmux_6_3_26866_26898 (
    .I(net_26866),
    .O(net_26898)
  );
  InMux inmux_6_3_26867_26900 (
    .I(net_26867),
    .O(net_26900)
  );
  ClkMux inmux_6_3_5_26896 (
    .I(net_5),
    .O(net_26896)
  );
  InMux inmux_6_4_26939_26991 (
    .I(net_26939),
    .O(net_26991)
  );
  InMux inmux_6_4_26943_27002 (
    .I(net_26943),
    .O(net_27002)
  );
  InMux inmux_6_4_26944_27007 (
    .I(net_26944),
    .O(net_27007)
  );
  InMux inmux_6_4_26945_27006 (
    .I(net_26945),
    .O(net_27006)
  );
  InMux inmux_6_4_26949_27005 (
    .I(net_26949),
    .O(net_27005)
  );
  CEMux inmux_6_4_26950_26999 (
    .I(net_26950),
    .O(net_26999)
  );
  InMux inmux_6_4_26951_27003 (
    .I(net_26951),
    .O(net_27003)
  );
  SRMux inmux_6_4_26952_27008 (
    .I(net_26952),
    .O(net_27008)
  );
  InMux inmux_6_4_26955_27000 (
    .I(net_26955),
    .O(net_27000)
  );
  InMux inmux_6_4_26956_26987 (
    .I(net_26956),
    .O(net_26987)
  );
  InMux inmux_6_4_26957_26979 (
    .I(net_26957),
    .O(net_26979)
  );
  InMux inmux_6_4_26957_26981 (
    .I(net_26957),
    .O(net_26981)
  );
  InMux inmux_6_4_26957_26983 (
    .I(net_26957),
    .O(net_26983)
  );
  InMux inmux_6_4_26957_26985 (
    .I(net_26957),
    .O(net_26985)
  );
  InMux inmux_6_4_26960_26992 (
    .I(net_26960),
    .O(net_26992)
  );
  InMux inmux_6_4_26961_26993 (
    .I(net_26961),
    .O(net_26993)
  );
  InMux inmux_6_4_26962_26990 (
    .I(net_26962),
    .O(net_26990)
  );
  InMux inmux_6_4_26964_27004 (
    .I(net_26964),
    .O(net_27004)
  );
  InMux inmux_6_4_26965_26980 (
    .I(net_26965),
    .O(net_26980)
  );
  InMux inmux_6_4_26965_26982 (
    .I(net_26965),
    .O(net_26982)
  );
  InMux inmux_6_4_26965_26984 (
    .I(net_26965),
    .O(net_26984)
  );
  InMux inmux_6_4_26965_26986 (
    .I(net_26965),
    .O(net_26986)
  );
  InMux inmux_6_4_26968_26988 (
    .I(net_26968),
    .O(net_26988)
  );
  InMux inmux_6_4_26969_27001 (
    .I(net_26969),
    .O(net_27001)
  );
  ClkMux inmux_6_4_5_26998 (
    .I(net_5),
    .O(net_26998)
  );
  CEMux inmux_6_9_27467_27509 (
    .I(net_27467),
    .O(net_27509)
  );
  SRMux inmux_6_9_27469_27510 (
    .I(net_27469),
    .O(net_27510)
  );
  InMux inmux_6_9_27471_27498 (
    .I(net_27471),
    .O(net_27498)
  );
  InMux inmux_6_9_27477_27497 (
    .I(net_27477),
    .O(net_27497)
  );
  ClkMux inmux_6_9_5_27508 (
    .I(net_5),
    .O(net_27508)
  );
  IoInMux inmux_7_0_29752_29728 (
    .I(net_29752),
    .O(net_29728)
  );
  InMux inmux_7_10_30946_31001 (
    .I(net_30946),
    .O(net_31001)
  );
  InMux inmux_7_10_30950_30993 (
    .I(net_30950),
    .O(net_30993)
  );
  InMux inmux_7_10_30958_31018 (
    .I(net_30958),
    .O(net_31018)
  );
  InMux inmux_7_10_30959_30988 (
    .I(net_30959),
    .O(net_30988)
  );
  InMux inmux_7_10_30963_30983 (
    .I(net_30963),
    .O(net_30983)
  );
  InMux inmux_7_10_30967_30975 (
    .I(net_30967),
    .O(net_30975)
  );
  InMux inmux_7_10_30969_31011 (
    .I(net_30969),
    .O(net_31011)
  );
  ClkMux inmux_7_10_5_31022 (
    .I(net_5),
    .O(net_31022)
  );
  SRMux inmux_7_10_9_31023 (
    .I(net_9),
    .O(net_31023)
  );
  InMux inmux_7_11_31071_31100 (
    .I(net_31071),
    .O(net_31100)
  );
  InMux inmux_7_11_31076_31117 (
    .I(net_31076),
    .O(net_31117)
  );
  InMux inmux_7_11_31079_31140 (
    .I(net_31079),
    .O(net_31140)
  );
  InMux inmux_7_11_31084_31123 (
    .I(net_31084),
    .O(net_31123)
  );
  InMux inmux_7_11_31086_31128 (
    .I(net_31086),
    .O(net_31128)
  );
  InMux inmux_7_11_31087_31134 (
    .I(net_31087),
    .O(net_31134)
  );
  InMux inmux_7_11_31091_31104 (
    .I(net_31091),
    .O(net_31104)
  );
  InMux inmux_7_11_31095_31111 (
    .I(net_31095),
    .O(net_31111)
  );
  ClkMux inmux_7_11_5_31145 (
    .I(net_5),
    .O(net_31145)
  );
  SRMux inmux_7_11_9_31146 (
    .I(net_9),
    .O(net_31146)
  );
  InMux inmux_7_12_31189_31234 (
    .I(net_31189),
    .O(net_31234)
  );
  InMux inmux_7_12_31190_31235 (
    .I(net_31190),
    .O(net_31235)
  );
  InMux inmux_7_12_31191_31222 (
    .I(net_31191),
    .O(net_31222)
  );
  InMux inmux_7_12_31192_31240 (
    .I(net_31192),
    .O(net_31240)
  );
  InMux inmux_7_12_31195_31241 (
    .I(net_31195),
    .O(net_31241)
  );
  InMux inmux_7_12_31196_31258 (
    .I(net_31196),
    .O(net_31258)
  );
  InMux inmux_7_12_31197_31228 (
    .I(net_31197),
    .O(net_31228)
  );
  InMux inmux_7_12_31198_31253 (
    .I(net_31198),
    .O(net_31253)
  );
  InMux inmux_7_12_31199_31259 (
    .I(net_31199),
    .O(net_31259)
  );
  InMux inmux_7_12_31201_31247 (
    .I(net_31201),
    .O(net_31247)
  );
  InMux inmux_7_12_31203_31252 (
    .I(net_31203),
    .O(net_31252)
  );
  InMux inmux_7_12_31207_31246 (
    .I(net_31207),
    .O(net_31246)
  );
  InMux inmux_7_12_31214_31229 (
    .I(net_31214),
    .O(net_31229)
  );
  InMux inmux_7_12_31217_31223 (
    .I(net_31217),
    .O(net_31223)
  );
  InMux inmux_7_12_31220_31230 (
    .I(net_31220),
    .O(net_31230)
  );
  InMux inmux_7_12_31226_31236 (
    .I(net_31226),
    .O(net_31236)
  );
  InMux inmux_7_12_31232_31242 (
    .I(net_31232),
    .O(net_31242)
  );
  InMux inmux_7_12_31238_31248 (
    .I(net_31238),
    .O(net_31248)
  );
  InMux inmux_7_12_31244_31254 (
    .I(net_31244),
    .O(net_31254)
  );
  InMux inmux_7_12_31250_31260 (
    .I(net_31250),
    .O(net_31260)
  );
  InMux inmux_7_12_31256_31266 (
    .I(net_31256),
    .O(net_31266)
  );
  InMux inmux_7_13_31312_31386 (
    .I(net_31312),
    .O(net_31386)
  );
  InMux inmux_7_13_31313_31368 (
    .I(net_31313),
    .O(net_31368)
  );
  InMux inmux_7_13_31314_31364 (
    .I(net_31314),
    .O(net_31364)
  );
  InMux inmux_7_13_31315_31382 (
    .I(net_31315),
    .O(net_31382)
  );
  InMux inmux_7_13_31319_31376 (
    .I(net_31319),
    .O(net_31376)
  );
  InMux inmux_7_13_31322_31344 (
    .I(net_31322),
    .O(net_31344)
  );
  InMux inmux_7_13_31331_31356 (
    .I(net_31331),
    .O(net_31356)
  );
  InMux inmux_7_13_31340_31353 (
    .I(net_31340),
    .O(net_31353)
  );
  ClkMux inmux_7_13_5_31391 (
    .I(net_5),
    .O(net_31391)
  );
  SRMux inmux_7_13_9_31392 (
    .I(net_9),
    .O(net_31392)
  );
  InMux inmux_7_14_31444_31494 (
    .I(net_31444),
    .O(net_31494)
  );
  InMux inmux_7_14_31445_31505 (
    .I(net_31445),
    .O(net_31505)
  );
  InMux inmux_7_14_31448_31511 (
    .I(net_31448),
    .O(net_31511)
  );
  InMux inmux_7_14_31459_31486 (
    .I(net_31459),
    .O(net_31486)
  );
  ClkMux inmux_7_14_5_31514 (
    .I(net_5),
    .O(net_31514)
  );
  SRMux inmux_7_14_9_31515 (
    .I(net_9),
    .O(net_31515)
  );
  InMux inmux_7_15_31557_31628 (
    .I(net_31557),
    .O(net_31628)
  );
  InMux inmux_7_15_31558_31598 (
    .I(net_31558),
    .O(net_31598)
  );
  InMux inmux_7_15_31559_31614 (
    .I(net_31559),
    .O(net_31614)
  );
  InMux inmux_7_15_31561_31592 (
    .I(net_31561),
    .O(net_31592)
  );
  InMux inmux_7_15_31561_31597 (
    .I(net_31561),
    .O(net_31597)
  );
  InMux inmux_7_15_31561_31604 (
    .I(net_31561),
    .O(net_31604)
  );
  InMux inmux_7_15_31562_31596 (
    .I(net_31562),
    .O(net_31596)
  );
  InMux inmux_7_15_31563_31633 (
    .I(net_31563),
    .O(net_31633)
  );
  InMux inmux_7_15_31564_31634 (
    .I(net_31564),
    .O(net_31634)
  );
  InMux inmux_7_15_31565_31617 (
    .I(net_31565),
    .O(net_31617)
  );
  InMux inmux_7_15_31566_31602 (
    .I(net_31566),
    .O(net_31602)
  );
  InMux inmux_7_15_31567_31622 (
    .I(net_31567),
    .O(net_31622)
  );
  InMux inmux_7_15_31568_31599 (
    .I(net_31568),
    .O(net_31599)
  );
  InMux inmux_7_15_31569_31608 (
    .I(net_31569),
    .O(net_31608)
  );
  InMux inmux_7_15_31569_31615 (
    .I(net_31569),
    .O(net_31615)
  );
  InMux inmux_7_15_31569_31620 (
    .I(net_31569),
    .O(net_31620)
  );
  InMux inmux_7_15_31569_31632 (
    .I(net_31569),
    .O(net_31632)
  );
  InMux inmux_7_15_31570_31609 (
    .I(net_31570),
    .O(net_31609)
  );
  InMux inmux_7_15_31571_31603 (
    .I(net_31571),
    .O(net_31603)
  );
  InMux inmux_7_15_31572_31616 (
    .I(net_31572),
    .O(net_31616)
  );
  InMux inmux_7_15_31573_31590 (
    .I(net_31573),
    .O(net_31590)
  );
  InMux inmux_7_15_31574_31593 (
    .I(net_31574),
    .O(net_31593)
  );
  InMux inmux_7_15_31575_31611 (
    .I(net_31575),
    .O(net_31611)
  );
  InMux inmux_7_15_31577_31623 (
    .I(net_31577),
    .O(net_31623)
  );
  InMux inmux_7_15_31578_31591 (
    .I(net_31578),
    .O(net_31591)
  );
  InMux inmux_7_15_31582_31635 (
    .I(net_31582),
    .O(net_31635)
  );
  InMux inmux_7_15_31583_31610 (
    .I(net_31583),
    .O(net_31610)
  );
  CEMux inmux_7_15_31584_31636 (
    .I(net_31584),
    .O(net_31636)
  );
  InMux inmux_7_15_31585_31605 (
    .I(net_31585),
    .O(net_31605)
  );
  InMux inmux_7_15_31586_31621 (
    .I(net_31586),
    .O(net_31621)
  );
  ClkMux inmux_7_15_5_31637 (
    .I(net_5),
    .O(net_31637)
  );
  SRMux inmux_7_15_9_31638 (
    .I(net_9),
    .O(net_31638)
  );
  InMux inmux_7_16_31696_31756 (
    .I(net_31696),
    .O(net_31756)
  );
  InMux inmux_7_16_31699_31716 (
    .I(net_31699),
    .O(net_31716)
  );
  InMux inmux_7_16_31701_31731 (
    .I(net_31701),
    .O(net_31731)
  );
  InMux inmux_7_16_31709_31727 (
    .I(net_31709),
    .O(net_31727)
  );
  InMux inmux_7_16_31711_31737 (
    .I(net_31711),
    .O(net_31737)
  );
  ClkMux inmux_7_16_5_31760 (
    .I(net_5),
    .O(net_31760)
  );
  SRMux inmux_7_16_9_31761 (
    .I(net_9),
    .O(net_31761)
  );
  InMux inmux_7_17_31805_31843 (
    .I(net_31805),
    .O(net_31843)
  );
  InMux inmux_7_17_31806_31837 (
    .I(net_31806),
    .O(net_31837)
  );
  InMux inmux_7_17_31807_31838 (
    .I(net_31807),
    .O(net_31838)
  );
  InMux inmux_7_17_31808_31844 (
    .I(net_31808),
    .O(net_31844)
  );
  InMux inmux_7_17_31811_31873 (
    .I(net_31811),
    .O(net_31873)
  );
  InMux inmux_7_17_31812_31867 (
    .I(net_31812),
    .O(net_31867)
  );
  InMux inmux_7_17_31813_31868 (
    .I(net_31813),
    .O(net_31868)
  );
  InMux inmux_7_17_31814_31850 (
    .I(net_31814),
    .O(net_31850)
  );
  InMux inmux_7_17_31816_31862 (
    .I(net_31816),
    .O(net_31862)
  );
  InMux inmux_7_17_31817_31849 (
    .I(net_31817),
    .O(net_31849)
  );
  InMux inmux_7_17_31818_31855 (
    .I(net_31818),
    .O(net_31855)
  );
  InMux inmux_7_17_31824_31861 (
    .I(net_31824),
    .O(net_31861)
  );
  InMux inmux_7_17_31832_31874 (
    .I(net_31832),
    .O(net_31874)
  );
  InMux inmux_7_17_31833_31856 (
    .I(net_31833),
    .O(net_31856)
  );
  InMux inmux_7_17_31871_31881 (
    .I(net_31871),
    .O(net_31881)
  );
  ClkMux inmux_7_17_5_31883 (
    .I(net_5),
    .O(net_31883)
  );
  SRMux inmux_7_17_9_31884 (
    .I(net_9),
    .O(net_31884)
  );
  InMux inmux_7_18_31932_31995 (
    .I(net_31932),
    .O(net_31995)
  );
  InMux inmux_7_18_31934_31991 (
    .I(net_31934),
    .O(net_31991)
  );
  InMux inmux_7_18_31937_31961 (
    .I(net_31937),
    .O(net_31961)
  );
  InMux inmux_7_18_31939_31971 (
    .I(net_31939),
    .O(net_31971)
  );
  InMux inmux_7_18_31954_31979 (
    .I(net_31954),
    .O(net_31979)
  );
  InMux inmux_7_18_31956_31986 (
    .I(net_31956),
    .O(net_31986)
  );
  ClkMux inmux_7_18_5_32006 (
    .I(net_5),
    .O(net_32006)
  );
  SRMux inmux_7_18_9_32007 (
    .I(net_9),
    .O(net_32007)
  );
  InMux inmux_7_19_32065_32113 (
    .I(net_32065),
    .O(net_32113)
  );
  InMux inmux_7_19_32070_32119 (
    .I(net_32070),
    .O(net_32119)
  );
  InMux inmux_7_19_32072_32102 (
    .I(net_32072),
    .O(net_32102)
  );
  InMux inmux_7_19_32074_32084 (
    .I(net_32074),
    .O(net_32084)
  );
  ClkMux inmux_7_19_5_32129 (
    .I(net_5),
    .O(net_32129)
  );
  SRMux inmux_7_19_9_32130 (
    .I(net_9),
    .O(net_32130)
  );
  InMux inmux_7_1_29823_29834 (
    .I(net_29823),
    .O(net_29834)
  );
  ClkMux inmux_7_1_5_29875 (
    .I(net_5),
    .O(net_29875)
  );
  SRMux inmux_7_1_9_29876 (
    .I(net_9),
    .O(net_29876)
  );
  InMux inmux_7_2_29961_30018 (
    .I(net_29961),
    .O(net_30018)
  );
  InMux inmux_7_2_29980_30003 (
    .I(net_29980),
    .O(net_30003)
  );
  InMux inmux_7_2_29983_30010 (
    .I(net_29983),
    .O(net_30010)
  );
  ClkMux inmux_7_2_5_30038 (
    .I(net_5),
    .O(net_30038)
  );
  SRMux inmux_7_2_9_30039 (
    .I(net_9),
    .O(net_30039)
  );
  InMux inmux_7_3_30081_30116 (
    .I(net_30081),
    .O(net_30116)
  );
  InMux inmux_7_3_30091_30139 (
    .I(net_30091),
    .O(net_30139)
  );
  InMux inmux_7_3_30104_30132 (
    .I(net_30104),
    .O(net_30132)
  );
  InMux inmux_7_3_30112_30126 (
    .I(net_30112),
    .O(net_30126)
  );
  ClkMux inmux_7_3_5_30161 (
    .I(net_5),
    .O(net_30161)
  );
  SRMux inmux_7_3_9_30162 (
    .I(net_9),
    .O(net_30162)
  );
  InMux inmux_7_4_30208_30237 (
    .I(net_30208),
    .O(net_30237)
  );
  InMux inmux_7_4_30211_30281 (
    .I(net_30211),
    .O(net_30281)
  );
  InMux inmux_7_4_30221_30269 (
    .I(net_30221),
    .O(net_30269)
  );
  InMux inmux_7_4_30224_30244 (
    .I(net_30224),
    .O(net_30244)
  );
  InMux inmux_7_4_30225_30255 (
    .I(net_30225),
    .O(net_30255)
  );
  InMux inmux_7_4_30232_30252 (
    .I(net_30232),
    .O(net_30252)
  );
  InMux inmux_7_4_30235_30268 (
    .I(net_30235),
    .O(net_30268)
  );
  ClkMux inmux_7_4_5_30284 (
    .I(net_5),
    .O(net_30284)
  );
  SRMux inmux_7_4_9_30285 (
    .I(net_9),
    .O(net_30285)
  );
  InMux inmux_7_5_30329_30362 (
    .I(net_30329),
    .O(net_30362)
  );
  InMux inmux_7_5_30329_30393 (
    .I(net_30329),
    .O(net_30393)
  );
  InMux inmux_7_5_30333_30374 (
    .I(net_30333),
    .O(net_30374)
  );
  InMux inmux_7_5_30336_30386 (
    .I(net_30336),
    .O(net_30386)
  );
  InMux inmux_7_5_30337_30361 (
    .I(net_30337),
    .O(net_30361)
  );
  InMux inmux_7_5_30337_30368 (
    .I(net_30337),
    .O(net_30368)
  );
  InMux inmux_7_5_30337_30373 (
    .I(net_30337),
    .O(net_30373)
  );
  InMux inmux_7_5_30337_30380 (
    .I(net_30337),
    .O(net_30380)
  );
  InMux inmux_7_5_30337_30392 (
    .I(net_30337),
    .O(net_30392)
  );
  InMux inmux_7_5_30341_30385 (
    .I(net_30341),
    .O(net_30385)
  );
  InMux inmux_7_5_30342_30398 (
    .I(net_30342),
    .O(net_30398)
  );
  InMux inmux_7_5_30343_30396 (
    .I(net_30343),
    .O(net_30396)
  );
  InMux inmux_7_5_30346_30378 (
    .I(net_30346),
    .O(net_30378)
  );
  InMux inmux_7_5_30348_30397 (
    .I(net_30348),
    .O(net_30397)
  );
  InMux inmux_7_5_30350_30387 (
    .I(net_30350),
    .O(net_30387)
  );
  InMux inmux_7_5_30354_30403 (
    .I(net_30354),
    .O(net_30403)
  );
  InMux inmux_7_5_30355_30399 (
    .I(net_30355),
    .O(net_30399)
  );
  InMux inmux_7_5_30358_30367 (
    .I(net_30358),
    .O(net_30367)
  );
  InMux inmux_7_5_30359_30369 (
    .I(net_30359),
    .O(net_30369)
  );
  InMux inmux_7_5_30365_30375 (
    .I(net_30365),
    .O(net_30375)
  );
  InMux inmux_7_5_30371_30381 (
    .I(net_30371),
    .O(net_30381)
  );
  ClkMux inmux_7_5_5_30407 (
    .I(net_5),
    .O(net_30407)
  );
  CEMux inmux_7_5_8_30406 (
    .I(net_8),
    .O(net_30406)
  );
  InMux inmux_7_6_30453_30501 (
    .I(net_30453),
    .O(net_30501)
  );
  InMux inmux_7_6_30455_30484 (
    .I(net_30455),
    .O(net_30484)
  );
  InMux inmux_7_6_30455_30525 (
    .I(net_30455),
    .O(net_30525)
  );
  InMux inmux_7_6_30459_30490 (
    .I(net_30459),
    .O(net_30490)
  );
  InMux inmux_7_6_30460_30496 (
    .I(net_30460),
    .O(net_30496)
  );
  InMux inmux_7_6_30461_30516 (
    .I(net_30461),
    .O(net_30516)
  );
  InMux inmux_7_6_30463_30485 (
    .I(net_30463),
    .O(net_30485)
  );
  InMux inmux_7_6_30463_30526 (
    .I(net_30463),
    .O(net_30526)
  );
  InMux inmux_7_6_30476_30508 (
    .I(net_30476),
    .O(net_30508)
  );
  InMux inmux_7_6_30477_30497 (
    .I(net_30477),
    .O(net_30497)
  );
  InMux inmux_7_6_30477_30502 (
    .I(net_30477),
    .O(net_30502)
  );
  InMux inmux_7_6_30478_30491 (
    .I(net_30478),
    .O(net_30491)
  );
  InMux inmux_7_6_30481_30521 (
    .I(net_30481),
    .O(net_30521)
  );
  InMux inmux_7_6_30482_30492 (
    .I(net_30482),
    .O(net_30492)
  );
  InMux inmux_7_6_30488_30498 (
    .I(net_30488),
    .O(net_30498)
  );
  InMux inmux_7_6_30494_30504 (
    .I(net_30494),
    .O(net_30504)
  );
  ClkMux inmux_7_6_5_30530 (
    .I(net_5),
    .O(net_30530)
  );
  SRMux inmux_7_6_9_30531 (
    .I(net_9),
    .O(net_30531)
  );
  InMux inmux_7_7_30575_30630 (
    .I(net_30575),
    .O(net_30630)
  );
  InMux inmux_7_7_30576_30636 (
    .I(net_30576),
    .O(net_30636)
  );
  InMux inmux_7_7_30579_30632 (
    .I(net_30579),
    .O(net_30632)
  );
  InMux inmux_7_7_30579_30639 (
    .I(net_30579),
    .O(net_30639)
  );
  InMux inmux_7_7_30580_30645 (
    .I(net_30580),
    .O(net_30645)
  );
  InMux inmux_7_7_30584_30608 (
    .I(net_30584),
    .O(net_30608)
  );
  InMux inmux_7_7_30591_30625 (
    .I(net_30591),
    .O(net_30625)
  );
  InMux inmux_7_7_30592_30614 (
    .I(net_30592),
    .O(net_30614)
  );
  InMux inmux_7_7_30601_30621 (
    .I(net_30601),
    .O(net_30621)
  );
  InMux inmux_7_7_30604_30649 (
    .I(net_30604),
    .O(net_30649)
  );
  ClkMux inmux_7_7_5_30653 (
    .I(net_5),
    .O(net_30653)
  );
  SRMux inmux_7_7_9_30654 (
    .I(net_9),
    .O(net_30654)
  );
  InMux inmux_7_8_30696_30760 (
    .I(net_30696),
    .O(net_30760)
  );
  InMux inmux_7_8_30702_30774 (
    .I(net_30702),
    .O(net_30774)
  );
  InMux inmux_7_8_30704_30735 (
    .I(net_30704),
    .O(net_30735)
  );
  InMux inmux_7_8_30712_30743 (
    .I(net_30712),
    .O(net_30743)
  );
  InMux inmux_7_8_30718_30755 (
    .I(net_30718),
    .O(net_30755)
  );
  InMux inmux_7_8_30720_30747 (
    .I(net_30720),
    .O(net_30747)
  );
  InMux inmux_7_8_30724_30732 (
    .I(net_30724),
    .O(net_30732)
  );
  InMux inmux_7_8_30726_30766 (
    .I(net_30726),
    .O(net_30766)
  );
  ClkMux inmux_7_8_5_30776 (
    .I(net_5),
    .O(net_30776)
  );
  SRMux inmux_7_8_9_30777 (
    .I(net_9),
    .O(net_30777)
  );
  CEMux inmux_7_9_10_30898 (
    .I(net_10),
    .O(net_30898)
  );
  InMux inmux_7_9_30820_30865 (
    .I(net_30820),
    .O(net_30865)
  );
  InMux inmux_7_9_30828_30852 (
    .I(net_30828),
    .O(net_30852)
  );
  InMux inmux_7_9_30830_30861 (
    .I(net_30830),
    .O(net_30861)
  );
  InMux inmux_7_9_30831_30896 (
    .I(net_30831),
    .O(net_30896)
  );
  InMux inmux_7_9_30836_30891 (
    .I(net_30836),
    .O(net_30891)
  );
  InMux inmux_7_9_30841_30873 (
    .I(net_30841),
    .O(net_30873)
  );
  InMux inmux_7_9_30848_30876 (
    .I(net_30848),
    .O(net_30876)
  );
  ClkMux inmux_7_9_5_30899 (
    .I(net_5),
    .O(net_30899)
  );
  IoInMux inmux_8_0_33572_33559 (
    .I(net_33572),
    .O(net_33559)
  );
  InMux inmux_8_10_34773_34813 (
    .I(net_34773),
    .O(net_34813)
  );
  InMux inmux_8_10_34788_34820 (
    .I(net_34788),
    .O(net_34820)
  );
  CEMux inmux_8_10_34791_34852 (
    .I(net_34791),
    .O(net_34852)
  );
  ClkMux inmux_8_10_5_34853 (
    .I(net_5),
    .O(net_34853)
  );
  InMux inmux_8_11_34904_34937 (
    .I(net_34904),
    .O(net_34937)
  );
  InMux inmux_8_11_34906_34968 (
    .I(net_34906),
    .O(net_34968)
  );
  InMux inmux_8_11_34908_34932 (
    .I(net_34908),
    .O(net_34932)
  );
  InMux inmux_8_11_34916_34953 (
    .I(net_34916),
    .O(net_34953)
  );
  InMux inmux_8_11_34918_34962 (
    .I(net_34918),
    .O(net_34962)
  );
  InMux inmux_8_11_34920_34947 (
    .I(net_34920),
    .O(net_34947)
  );
  InMux inmux_8_11_34922_34971 (
    .I(net_34922),
    .O(net_34971)
  );
  InMux inmux_8_11_34926_34942 (
    .I(net_34926),
    .O(net_34942)
  );
  ClkMux inmux_8_11_5_34976 (
    .I(net_5),
    .O(net_34976)
  );
  SRMux inmux_8_11_9_34977 (
    .I(net_9),
    .O(net_34977)
  );
  InMux inmux_8_12_35021_35066 (
    .I(net_35021),
    .O(net_35066)
  );
  InMux inmux_8_12_35023_35078 (
    .I(net_35023),
    .O(net_35078)
  );
  InMux inmux_8_12_35028_35059 (
    .I(net_35028),
    .O(net_35059)
  );
  InMux inmux_8_12_35030_35071 (
    .I(net_35030),
    .O(net_35071)
  );
  InMux inmux_8_12_35032_35083 (
    .I(net_35032),
    .O(net_35083)
  );
  InMux inmux_8_12_35033_35089 (
    .I(net_35033),
    .O(net_35089)
  );
  InMux inmux_8_12_35034_35095 (
    .I(net_35034),
    .O(net_35095)
  );
  InMux inmux_8_12_35035_35054 (
    .I(net_35035),
    .O(net_35054)
  );
  InMux inmux_8_12_35040_35053 (
    .I(net_35040),
    .O(net_35053)
  );
  InMux inmux_8_12_35087_35097 (
    .I(net_35087),
    .O(net_35097)
  );
  ClkMux inmux_8_12_5_35099 (
    .I(net_5),
    .O(net_35099)
  );
  SRMux inmux_8_12_9_35100 (
    .I(net_9),
    .O(net_35100)
  );
  InMux inmux_8_13_35137_35178 (
    .I(net_35137),
    .O(net_35178)
  );
  InMux inmux_8_13_35154_35207 (
    .I(net_35154),
    .O(net_35207)
  );
  InMux inmux_8_13_35158_35218 (
    .I(net_35158),
    .O(net_35218)
  );
  InMux inmux_8_13_35161_35202 (
    .I(net_35161),
    .O(net_35202)
  );
  InMux inmux_8_13_35168_35212 (
    .I(net_35168),
    .O(net_35212)
  );
  InMux inmux_8_13_35170_35181 (
    .I(net_35170),
    .O(net_35181)
  );
  InMux inmux_8_13_35172_35193 (
    .I(net_35172),
    .O(net_35193)
  );
  InMux inmux_8_13_35173_35189 (
    .I(net_35173),
    .O(net_35189)
  );
  ClkMux inmux_8_13_5_35222 (
    .I(net_5),
    .O(net_35222)
  );
  SRMux inmux_8_13_9_35223 (
    .I(net_9),
    .O(net_35223)
  );
  InMux inmux_8_14_35269_35298 (
    .I(net_35269),
    .O(net_35298)
  );
  InMux inmux_8_14_35273_35337 (
    .I(net_35273),
    .O(net_35337)
  );
  InMux inmux_8_14_35276_35334 (
    .I(net_35276),
    .O(net_35334)
  );
  InMux inmux_8_14_35281_35336 (
    .I(net_35281),
    .O(net_35336)
  );
  InMux inmux_8_14_35282_35335 (
    .I(net_35282),
    .O(net_35335)
  );
  ClkMux inmux_8_14_5_35345 (
    .I(net_5),
    .O(net_35345)
  );
  CEMux inmux_8_14_8_35344 (
    .I(net_8),
    .O(net_35344)
  );
  InMux inmux_8_15_35388_35428 (
    .I(net_35388),
    .O(net_35428)
  );
  InMux inmux_8_15_35390_35440 (
    .I(net_35390),
    .O(net_35440)
  );
  InMux inmux_8_15_35391_35460 (
    .I(net_35391),
    .O(net_35460)
  );
  InMux inmux_8_15_35392_35445 (
    .I(net_35392),
    .O(net_35445)
  );
  InMux inmux_8_15_35394_35423 (
    .I(net_35394),
    .O(net_35423)
  );
  InMux inmux_8_15_35396_35441 (
    .I(net_35396),
    .O(net_35441)
  );
  InMux inmux_8_15_35397_35442 (
    .I(net_35397),
    .O(net_35442)
  );
  InMux inmux_8_15_35399_35457 (
    .I(net_35399),
    .O(net_35457)
  );
  InMux inmux_8_15_35400_35422 (
    .I(net_35400),
    .O(net_35422)
  );
  InMux inmux_8_15_35401_35466 (
    .I(net_35401),
    .O(net_35466)
  );
  InMux inmux_8_15_35402_35434 (
    .I(net_35402),
    .O(net_35434)
  );
  InMux inmux_8_15_35403_35430 (
    .I(net_35403),
    .O(net_35430)
  );
  InMux inmux_8_15_35404_35421 (
    .I(net_35404),
    .O(net_35421)
  );
  InMux inmux_8_15_35405_35446 (
    .I(net_35405),
    .O(net_35446)
  );
  CEMux inmux_8_15_35406_35467 (
    .I(net_35406),
    .O(net_35467)
  );
  InMux inmux_8_15_35407_35424 (
    .I(net_35407),
    .O(net_35424)
  );
  InMux inmux_8_15_35407_35427 (
    .I(net_35407),
    .O(net_35427)
  );
  InMux inmux_8_15_35407_35436 (
    .I(net_35407),
    .O(net_35436)
  );
  InMux inmux_8_15_35407_35439 (
    .I(net_35407),
    .O(net_35439)
  );
  InMux inmux_8_15_35407_35448 (
    .I(net_35407),
    .O(net_35448)
  );
  InMux inmux_8_15_35407_35458 (
    .I(net_35407),
    .O(net_35458)
  );
  InMux inmux_8_15_35407_35465 (
    .I(net_35407),
    .O(net_35465)
  );
  InMux inmux_8_15_35410_35459 (
    .I(net_35410),
    .O(net_35459)
  );
  InMux inmux_8_15_35413_35433 (
    .I(net_35413),
    .O(net_35433)
  );
  InMux inmux_8_15_35414_35429 (
    .I(net_35414),
    .O(net_35429)
  );
  InMux inmux_8_15_35415_35447 (
    .I(net_35415),
    .O(net_35447)
  );
  InMux inmux_8_15_35416_35463 (
    .I(net_35416),
    .O(net_35463)
  );
  InMux inmux_8_15_35417_35464 (
    .I(net_35417),
    .O(net_35464)
  );
  InMux inmux_8_15_35419_35435 (
    .I(net_35419),
    .O(net_35435)
  );
  ClkMux inmux_8_15_5_35468 (
    .I(net_5),
    .O(net_35468)
  );
  InMux inmux_8_16_35513_35565 (
    .I(net_35513),
    .O(net_35565)
  );
  InMux inmux_8_16_35515_35551 (
    .I(net_35515),
    .O(net_35551)
  );
  InMux inmux_8_16_35519_35581 (
    .I(net_35519),
    .O(net_35581)
  );
  CEMux inmux_8_16_35522_35590 (
    .I(net_35522),
    .O(net_35590)
  );
  InMux inmux_8_16_35524_35580 (
    .I(net_35524),
    .O(net_35580)
  );
  InMux inmux_8_16_35525_35552 (
    .I(net_35525),
    .O(net_35552)
  );
  InMux inmux_8_16_35526_35582 (
    .I(net_35526),
    .O(net_35582)
  );
  InMux inmux_8_16_35528_35564 (
    .I(net_35528),
    .O(net_35564)
  );
  InMux inmux_8_16_35528_35583 (
    .I(net_35528),
    .O(net_35583)
  );
  InMux inmux_8_16_35530_35550 (
    .I(net_35530),
    .O(net_35550)
  );
  InMux inmux_8_16_35533_35563 (
    .I(net_35533),
    .O(net_35563)
  );
  InMux inmux_8_16_35535_35562 (
    .I(net_35535),
    .O(net_35562)
  );
  InMux inmux_8_16_35536_35553 (
    .I(net_35536),
    .O(net_35553)
  );
  ClkMux inmux_8_16_5_35591 (
    .I(net_5),
    .O(net_35591)
  );
  SRMux inmux_8_16_9_35592 (
    .I(net_9),
    .O(net_35592)
  );
  InMux inmux_8_1_33635_33695 (
    .I(net_33635),
    .O(net_33695)
  );
  InMux inmux_8_1_33644_33678 (
    .I(net_33644),
    .O(net_33678)
  );
  InMux inmux_8_1_33646_33673 (
    .I(net_33646),
    .O(net_33673)
  );
  InMux inmux_8_1_33648_33704 (
    .I(net_33648),
    .O(net_33704)
  );
  InMux inmux_8_1_33652_33689 (
    .I(net_33652),
    .O(net_33689)
  );
  ClkMux inmux_8_1_5_33706 (
    .I(net_5),
    .O(net_33706)
  );
  SRMux inmux_8_1_9_33707 (
    .I(net_9),
    .O(net_33707)
  );
  InMux inmux_8_2_33812_33835 (
    .I(net_33812),
    .O(net_33835)
  );
  InMux inmux_8_2_33813_33859 (
    .I(net_33813),
    .O(net_33859)
  );
  InMux inmux_8_2_33818_33824 (
    .I(net_33818),
    .O(net_33824)
  );
  ClkMux inmux_8_2_5_33869 (
    .I(net_5),
    .O(net_33869)
  );
  SRMux inmux_8_2_9_33870 (
    .I(net_9),
    .O(net_33870)
  );
  CEMux inmux_8_3_33914_33991 (
    .I(net_33914),
    .O(net_33991)
  );
  InMux inmux_8_3_33917_33982 (
    .I(net_33917),
    .O(net_33982)
  );
  InMux inmux_8_3_33918_33945 (
    .I(net_33918),
    .O(net_33945)
  );
  InMux inmux_8_3_33931_33946 (
    .I(net_33931),
    .O(net_33946)
  );
  InMux inmux_8_3_33931_33984 (
    .I(net_33931),
    .O(net_33984)
  );
  InMux inmux_8_3_33933_33975 (
    .I(net_33933),
    .O(net_33975)
  );
  InMux inmux_8_3_33934_33981 (
    .I(net_33934),
    .O(net_33981)
  );
  InMux inmux_8_3_33935_33948 (
    .I(net_33935),
    .O(net_33948)
  );
  InMux inmux_8_3_33937_33947 (
    .I(net_33937),
    .O(net_33947)
  );
  InMux inmux_8_3_33937_33983 (
    .I(net_33937),
    .O(net_33983)
  );
  InMux inmux_8_3_33941_33990 (
    .I(net_33941),
    .O(net_33990)
  );
  ClkMux inmux_8_3_5_33992 (
    .I(net_5),
    .O(net_33992)
  );
  InMux inmux_8_4_34038_34086 (
    .I(net_34038),
    .O(net_34086)
  );
  InMux inmux_8_4_34040_34071 (
    .I(net_34040),
    .O(net_34071)
  );
  InMux inmux_8_4_34045_34107 (
    .I(net_34045),
    .O(net_34107)
  );
  InMux inmux_8_4_34053_34099 (
    .I(net_34053),
    .O(net_34099)
  );
  InMux inmux_8_4_34055_34092 (
    .I(net_34055),
    .O(net_34092)
  );
  InMux inmux_8_4_34056_34110 (
    .I(net_34056),
    .O(net_34110)
  );
  InMux inmux_8_4_34064_34080 (
    .I(net_34064),
    .O(net_34080)
  );
  ClkMux inmux_8_4_5_34115 (
    .I(net_5),
    .O(net_34115)
  );
  SRMux inmux_8_4_9_34116 (
    .I(net_9),
    .O(net_34116)
  );
  InMux inmux_8_5_34160_34227 (
    .I(net_34160),
    .O(net_34227)
  );
  InMux inmux_8_5_34167_34205 (
    .I(net_34167),
    .O(net_34205)
  );
  InMux inmux_8_5_34171_34215 (
    .I(net_34171),
    .O(net_34215)
  );
  InMux inmux_8_5_34171_34222 (
    .I(net_34171),
    .O(net_34222)
  );
  InMux inmux_8_5_34179_34192 (
    .I(net_34179),
    .O(net_34192)
  );
  InMux inmux_8_5_34181_34197 (
    .I(net_34181),
    .O(net_34197)
  );
  InMux inmux_8_5_34185_34217 (
    .I(net_34185),
    .O(net_34217)
  );
  InMux inmux_8_5_34186_34235 (
    .I(net_34186),
    .O(net_34235)
  );
  InMux inmux_8_5_34187_34212 (
    .I(net_34187),
    .O(net_34212)
  );
  InMux inmux_8_5_34189_34224 (
    .I(net_34189),
    .O(net_34224)
  );
  ClkMux inmux_8_5_5_34238 (
    .I(net_5),
    .O(net_34238)
  );
  SRMux inmux_8_5_9_34239 (
    .I(net_9),
    .O(net_34239)
  );
  CEMux inmux_8_6_12_34360 (
    .I(net_12),
    .O(net_34360)
  );
  InMux inmux_8_6_34284_34332 (
    .I(net_34284),
    .O(net_34332)
  );
  InMux inmux_8_6_34286_34346 (
    .I(net_34286),
    .O(net_34346)
  );
  InMux inmux_8_6_34294_34314 (
    .I(net_34294),
    .O(net_34314)
  );
  InMux inmux_8_6_34298_34356 (
    .I(net_34298),
    .O(net_34356)
  );
  InMux inmux_8_6_34300_34353 (
    .I(net_34300),
    .O(net_34353)
  );
  InMux inmux_8_6_34304_34341 (
    .I(net_34304),
    .O(net_34341)
  );
  InMux inmux_8_6_34306_34323 (
    .I(net_34306),
    .O(net_34323)
  );
  ClkMux inmux_8_6_5_34361 (
    .I(net_5),
    .O(net_34361)
  );
  CEMux inmux_8_7_10_34483 (
    .I(net_10),
    .O(net_34483)
  );
  InMux inmux_8_7_34406_34439 (
    .I(net_34406),
    .O(net_34439)
  );
  InMux inmux_8_7_34409_34476 (
    .I(net_34409),
    .O(net_34476)
  );
  InMux inmux_8_7_34418_34450 (
    .I(net_34418),
    .O(net_34450)
  );
  ClkMux inmux_8_7_5_34484 (
    .I(net_5),
    .O(net_34484)
  );
  InMux inmux_8_8_34528_34573 (
    .I(net_34528),
    .O(net_34573)
  );
  InMux inmux_8_8_34529_34586 (
    .I(net_34529),
    .O(net_34586)
  );
  InMux inmux_8_8_34531_34579 (
    .I(net_34531),
    .O(net_34579)
  );
  InMux inmux_8_8_34532_34597 (
    .I(net_34532),
    .O(net_34597)
  );
  InMux inmux_8_8_34534_34592 (
    .I(net_34534),
    .O(net_34592)
  );
  InMux inmux_8_8_34539_34561 (
    .I(net_34539),
    .O(net_34561)
  );
  InMux inmux_8_8_34540_34574 (
    .I(net_34540),
    .O(net_34574)
  );
  InMux inmux_8_8_34541_34585 (
    .I(net_34541),
    .O(net_34585)
  );
  InMux inmux_8_8_34542_34562 (
    .I(net_34542),
    .O(net_34562)
  );
  InMux inmux_8_8_34544_34568 (
    .I(net_34544),
    .O(net_34568)
  );
  InMux inmux_8_8_34547_34598 (
    .I(net_34547),
    .O(net_34598)
  );
  InMux inmux_8_8_34552_34567 (
    .I(net_34552),
    .O(net_34567)
  );
  InMux inmux_8_8_34553_34580 (
    .I(net_34553),
    .O(net_34580)
  );
  InMux inmux_8_8_34558_34591 (
    .I(net_34558),
    .O(net_34591)
  );
  InMux inmux_8_8_34559_34569 (
    .I(net_34559),
    .O(net_34569)
  );
  InMux inmux_8_8_34565_34575 (
    .I(net_34565),
    .O(net_34575)
  );
  InMux inmux_8_8_34571_34581 (
    .I(net_34571),
    .O(net_34581)
  );
  InMux inmux_8_8_34577_34587 (
    .I(net_34577),
    .O(net_34587)
  );
  InMux inmux_8_8_34583_34593 (
    .I(net_34583),
    .O(net_34593)
  );
  InMux inmux_8_8_34589_34599 (
    .I(net_34589),
    .O(net_34599)
  );
  InMux inmux_8_8_34595_34605 (
    .I(net_34595),
    .O(net_34605)
  );
  InMux inmux_8_9_34652_34726 (
    .I(net_34652),
    .O(net_34726)
  );
  InMux inmux_8_9_34662_34691 (
    .I(net_34662),
    .O(net_34691)
  );
  InMux inmux_8_9_34664_34696 (
    .I(net_34664),
    .O(net_34696)
  );
  InMux inmux_8_9_34665_34692 (
    .I(net_34665),
    .O(net_34692)
  );
  InMux inmux_8_9_34668_34714 (
    .I(net_34668),
    .O(net_34714)
  );
  InMux inmux_8_9_34672_34709 (
    .I(net_34672),
    .O(net_34709)
  );
  InMux inmux_8_9_34676_34686 (
    .I(net_34676),
    .O(net_34686)
  );
  InMux inmux_8_9_34678_34722 (
    .I(net_34678),
    .O(net_34722)
  );
  ClkMux inmux_8_9_5_34730 (
    .I(net_5),
    .O(net_34730)
  );
  SRMux inmux_8_9_9_34731 (
    .I(net_9),
    .O(net_34731)
  );
  IoInMux inmux_9_0_37403_37390 (
    .I(net_37403),
    .O(net_37390)
  );
  IoInMux inmux_9_0_37406_37393 (
    .I(net_37406),
    .O(net_37393)
  );
  InMux inmux_9_10_38604_38649 (
    .I(net_38604),
    .O(net_38649)
  );
  InMux inmux_9_10_38608_38670 (
    .I(net_38608),
    .O(net_38670)
  );
  InMux inmux_9_10_38614_38662 (
    .I(net_38614),
    .O(net_38662)
  );
  InMux inmux_9_10_38615_38675 (
    .I(net_38615),
    .O(net_38675)
  );
  InMux inmux_9_10_38616_38679 (
    .I(net_38616),
    .O(net_38679)
  );
  InMux inmux_9_10_38624_38639 (
    .I(net_38624),
    .O(net_38639)
  );
  InMux inmux_9_10_38629_38680 (
    .I(net_38629),
    .O(net_38680)
  );
  InMux inmux_9_10_38632_38643 (
    .I(net_38632),
    .O(net_38643)
  );
  ClkMux inmux_9_10_5_38684 (
    .I(net_5),
    .O(net_38684)
  );
  SRMux inmux_9_10_9_38685 (
    .I(net_9),
    .O(net_38685)
  );
  InMux inmux_9_11_38735_38761 (
    .I(net_38735),
    .O(net_38761)
  );
  InMux inmux_9_11_38735_38797 (
    .I(net_38735),
    .O(net_38797)
  );
  CEMux inmux_9_11_38738_38806 (
    .I(net_38738),
    .O(net_38806)
  );
  InMux inmux_9_11_38749_38760 (
    .I(net_38749),
    .O(net_38760)
  );
  InMux inmux_9_11_38749_38796 (
    .I(net_38749),
    .O(net_38796)
  );
  ClkMux inmux_9_11_5_38807 (
    .I(net_5),
    .O(net_38807)
  );
  SRMux inmux_9_11_9_38808 (
    .I(net_9),
    .O(net_38808)
  );
  CEMux inmux_9_12_38852_38929 (
    .I(net_38852),
    .O(net_38929)
  );
  InMux inmux_9_12_38858_38891 (
    .I(net_38858),
    .O(net_38891)
  );
  InMux inmux_9_12_38873_38886 (
    .I(net_38873),
    .O(net_38886)
  );
  InMux inmux_9_12_38877_38916 (
    .I(net_38877),
    .O(net_38916)
  );
  InMux inmux_9_12_38879_38914 (
    .I(net_38879),
    .O(net_38914)
  );
  InMux inmux_9_12_38880_38908 (
    .I(net_38880),
    .O(net_38908)
  );
  ClkMux inmux_9_12_5_38930 (
    .I(net_5),
    .O(net_38930)
  );
  InMux inmux_9_13_38982_39042 (
    .I(net_38982),
    .O(net_39042)
  );
  InMux inmux_9_13_38983_39026 (
    .I(net_38983),
    .O(net_39026)
  );
  InMux inmux_9_13_38984_39039 (
    .I(net_38984),
    .O(net_39039)
  );
  InMux inmux_9_13_38990_39043 (
    .I(net_38990),
    .O(net_39043)
  );
  CEMux inmux_9_13_38991_39052 (
    .I(net_38991),
    .O(net_39052)
  );
  InMux inmux_9_13_39000_39044 (
    .I(net_39000),
    .O(net_39044)
  );
  InMux inmux_9_13_39003_39045 (
    .I(net_39003),
    .O(net_39045)
  );
  ClkMux inmux_9_13_5_39053 (
    .I(net_5),
    .O(net_39053)
  );
  InMux inmux_9_14_39098_39131 (
    .I(net_39098),
    .O(net_39131)
  );
  InMux inmux_9_14_39099_39156 (
    .I(net_39099),
    .O(net_39156)
  );
  InMux inmux_9_14_39100_39129 (
    .I(net_39100),
    .O(net_39129)
  );
  InMux inmux_9_14_39107_39148 (
    .I(net_39107),
    .O(net_39148)
  );
  InMux inmux_9_14_39110_39171 (
    .I(net_39110),
    .O(net_39171)
  );
  InMux inmux_9_14_39114_39162 (
    .I(net_39114),
    .O(net_39162)
  );
  InMux inmux_9_14_39115_39132 (
    .I(net_39115),
    .O(net_39132)
  );
  InMux inmux_9_14_39118_39141 (
    .I(net_39118),
    .O(net_39141)
  );
  CEMux inmux_9_14_39123_39175 (
    .I(net_39123),
    .O(net_39175)
  );
  InMux inmux_9_14_39126_39130 (
    .I(net_39126),
    .O(net_39130)
  );
  ClkMux inmux_9_14_5_39176 (
    .I(net_5),
    .O(net_39176)
  );
  InMux inmux_9_15_39224_39294 (
    .I(net_39224),
    .O(net_39294)
  );
  InMux inmux_9_15_39228_39254 (
    .I(net_39228),
    .O(net_39254)
  );
  CEMux inmux_9_15_39230_39298 (
    .I(net_39230),
    .O(net_39298)
  );
  InMux inmux_9_15_39231_39277 (
    .I(net_39231),
    .O(net_39277)
  );
  InMux inmux_9_15_39233_39260 (
    .I(net_39233),
    .O(net_39260)
  );
  InMux inmux_9_15_39233_39279 (
    .I(net_39233),
    .O(net_39279)
  );
  InMux inmux_9_15_39234_39261 (
    .I(net_39234),
    .O(net_39261)
  );
  InMux inmux_9_15_39235_39276 (
    .I(net_39235),
    .O(net_39276)
  );
  InMux inmux_9_15_39236_39291 (
    .I(net_39236),
    .O(net_39291)
  );
  InMux inmux_9_15_39238_39284 (
    .I(net_39238),
    .O(net_39284)
  );
  InMux inmux_9_15_39244_39259 (
    .I(net_39244),
    .O(net_39259)
  );
  InMux inmux_9_15_39244_39278 (
    .I(net_39244),
    .O(net_39278)
  );
  InMux inmux_9_15_39246_39266 (
    .I(net_39246),
    .O(net_39266)
  );
  InMux inmux_9_15_39247_39258 (
    .I(net_39247),
    .O(net_39258)
  );
  InMux inmux_9_15_39249_39272 (
    .I(net_39249),
    .O(net_39272)
  );
  ClkMux inmux_9_15_5_39299 (
    .I(net_5),
    .O(net_39299)
  );
  CEMux inmux_9_16_39344_39421 (
    .I(net_39344),
    .O(net_39421)
  );
  InMux inmux_9_16_39345_39376 (
    .I(net_39345),
    .O(net_39376)
  );
  InMux inmux_9_16_39348_39394 (
    .I(net_39348),
    .O(net_39394)
  );
  InMux inmux_9_16_39352_39419 (
    .I(net_39352),
    .O(net_39419)
  );
  InMux inmux_9_16_39360_39406 (
    .I(net_39360),
    .O(net_39406)
  );
  InMux inmux_9_16_39364_39401 (
    .I(net_39364),
    .O(net_39401)
  );
  ClkMux inmux_9_16_5_39422 (
    .I(net_5),
    .O(net_39422)
  );
  InMux inmux_9_17_39466_39506 (
    .I(net_39466),
    .O(net_39506)
  );
  InMux inmux_9_17_39466_39511 (
    .I(net_39466),
    .O(net_39511)
  );
  InMux inmux_9_17_39474_39507 (
    .I(net_39474),
    .O(net_39507)
  );
  InMux inmux_9_17_39476_39512 (
    .I(net_39476),
    .O(net_39512)
  );
  InMux inmux_9_17_39480_39498 (
    .I(net_39480),
    .O(net_39498)
  );
  InMux inmux_9_17_39481_39510 (
    .I(net_39481),
    .O(net_39510)
  );
  InMux inmux_9_17_39482_39518 (
    .I(net_39482),
    .O(net_39518)
  );
  CEMux inmux_9_17_39483_39544 (
    .I(net_39483),
    .O(net_39544)
  );
  InMux inmux_9_17_39484_39504 (
    .I(net_39484),
    .O(net_39504)
  );
  InMux inmux_9_17_39484_39513 (
    .I(net_39484),
    .O(net_39513)
  );
  InMux inmux_9_17_39492_39505 (
    .I(net_39492),
    .O(net_39505)
  );
  ClkMux inmux_9_17_5_39545 (
    .I(net_5),
    .O(net_39545)
  );
  InMux inmux_9_18_39588_39628 (
    .I(net_39588),
    .O(net_39628)
  );
  InMux inmux_9_18_39588_39635 (
    .I(net_39588),
    .O(net_39635)
  );
  InMux inmux_9_18_39589_39634 (
    .I(net_39589),
    .O(net_39634)
  );
  InMux inmux_9_18_39590_39623 (
    .I(net_39590),
    .O(net_39623)
  );
  InMux inmux_9_18_39591_39665 (
    .I(net_39591),
    .O(net_39665)
  );
  InMux inmux_9_18_39592_39657 (
    .I(net_39592),
    .O(net_39657)
  );
  InMux inmux_9_18_39594_39654 (
    .I(net_39594),
    .O(net_39654)
  );
  InMux inmux_9_18_39595_39627 (
    .I(net_39595),
    .O(net_39627)
  );
  InMux inmux_9_18_39596_39629 (
    .I(net_39596),
    .O(net_39629)
  );
  InMux inmux_9_18_39597_39664 (
    .I(net_39597),
    .O(net_39664)
  );
  InMux inmux_9_18_39598_39658 (
    .I(net_39598),
    .O(net_39658)
  );
  CEMux inmux_9_18_39599_39667 (
    .I(net_39599),
    .O(net_39667)
  );
  InMux inmux_9_18_39600_39622 (
    .I(net_39600),
    .O(net_39622)
  );
  InMux inmux_9_18_39602_39636 (
    .I(net_39602),
    .O(net_39636)
  );
  InMux inmux_9_18_39603_39630 (
    .I(net_39603),
    .O(net_39630)
  );
  InMux inmux_9_18_39604_39633 (
    .I(net_39604),
    .O(net_39633)
  );
  InMux inmux_9_18_39608_39666 (
    .I(net_39608),
    .O(net_39666)
  );
  InMux inmux_9_18_39610_39652 (
    .I(net_39610),
    .O(net_39652)
  );
  InMux inmux_9_18_39612_39624 (
    .I(net_39612),
    .O(net_39624)
  );
  InMux inmux_9_18_39612_39651 (
    .I(net_39612),
    .O(net_39651)
  );
  InMux inmux_9_18_39612_39660 (
    .I(net_39612),
    .O(net_39660)
  );
  InMux inmux_9_18_39612_39663 (
    .I(net_39612),
    .O(net_39663)
  );
  InMux inmux_9_18_39613_39621 (
    .I(net_39613),
    .O(net_39621)
  );
  InMux inmux_9_18_39615_39659 (
    .I(net_39615),
    .O(net_39659)
  );
  InMux inmux_9_18_39618_39653 (
    .I(net_39618),
    .O(net_39653)
  );
  ClkMux inmux_9_18_5_39668 (
    .I(net_5),
    .O(net_39668)
  );
  InMux inmux_9_1_37457_37533 (
    .I(net_37457),
    .O(net_37533)
  );
  InMux inmux_9_1_37462_37529 (
    .I(net_37462),
    .O(net_37529)
  );
  InMux inmux_9_1_37464_37498 (
    .I(net_37464),
    .O(net_37498)
  );
  InMux inmux_9_1_37468_37516 (
    .I(net_37468),
    .O(net_37516)
  );
  InMux inmux_9_1_37480_37510 (
    .I(net_37480),
    .O(net_37510)
  );
  ClkMux inmux_9_1_5_37537 (
    .I(net_5),
    .O(net_37537)
  );
  SRMux inmux_9_1_9_37538 (
    .I(net_9),
    .O(net_37538)
  );
  InMux inmux_9_2_37631_37672 (
    .I(net_37631),
    .O(net_37672)
  );
  InMux inmux_9_2_37633_37691 (
    .I(net_37633),
    .O(net_37691)
  );
  ClkMux inmux_9_2_5_37700 (
    .I(net_5),
    .O(net_37700)
  );
  CEMux inmux_9_2_8_37699 (
    .I(net_8),
    .O(net_37699)
  );
  InMux inmux_9_3_37743_37812 (
    .I(net_37743),
    .O(net_37812)
  );
  InMux inmux_9_3_37746_37815 (
    .I(net_37746),
    .O(net_37815)
  );
  InMux inmux_9_3_37749_37795 (
    .I(net_37749),
    .O(net_37795)
  );
  InMux inmux_9_3_37752_37814 (
    .I(net_37752),
    .O(net_37814)
  );
  CEMux inmux_9_3_37754_37822 (
    .I(net_37754),
    .O(net_37822)
  );
  InMux inmux_9_3_37762_37813 (
    .I(net_37762),
    .O(net_37813)
  );
  ClkMux inmux_9_3_5_37823 (
    .I(net_5),
    .O(net_37823)
  );
  CEMux inmux_9_4_37868_37945 (
    .I(net_37868),
    .O(net_37945)
  );
  InMux inmux_9_4_37870_37937 (
    .I(net_37870),
    .O(net_37937)
  );
  InMux inmux_9_4_37872_37942 (
    .I(net_37872),
    .O(net_37942)
  );
  InMux inmux_9_4_37873_37929 (
    .I(net_37873),
    .O(net_37929)
  );
  InMux inmux_9_4_37876_37914 (
    .I(net_37876),
    .O(net_37914)
  );
  InMux inmux_9_4_37880_37902 (
    .I(net_37880),
    .O(net_37902)
  );
  InMux inmux_9_4_37884_37899 (
    .I(net_37884),
    .O(net_37899)
  );
  InMux inmux_9_4_37885_37900 (
    .I(net_37885),
    .O(net_37900)
  );
  InMux inmux_9_4_37895_37901 (
    .I(net_37895),
    .O(net_37901)
  );
  ClkMux inmux_9_4_5_37946 (
    .I(net_5),
    .O(net_37946)
  );
  InMux inmux_9_5_37989_38041 (
    .I(net_37989),
    .O(net_38041)
  );
  InMux inmux_9_5_37989_38060 (
    .I(net_37989),
    .O(net_38060)
  );
  InMux inmux_9_5_37995_38058 (
    .I(net_37995),
    .O(net_38058)
  );
  InMux inmux_9_5_37997_38040 (
    .I(net_37997),
    .O(net_38040)
  );
  InMux inmux_9_5_37998_38024 (
    .I(net_37998),
    .O(net_38024)
  );
  InMux inmux_9_5_38008_38047 (
    .I(net_38008),
    .O(net_38047)
  );
  InMux inmux_9_5_38011_38031 (
    .I(net_38011),
    .O(net_38031)
  );
  InMux inmux_9_5_38016_38065 (
    .I(net_38016),
    .O(net_38065)
  );
  ClkMux inmux_9_5_5_38069 (
    .I(net_5),
    .O(net_38069)
  );
  SRMux inmux_9_5_9_38070 (
    .I(net_9),
    .O(net_38070)
  );
  InMux inmux_9_6_38118_38166 (
    .I(net_38118),
    .O(net_38166)
  );
  InMux inmux_9_6_38119_38160 (
    .I(net_38119),
    .O(net_38160)
  );
  InMux inmux_9_6_38120_38172 (
    .I(net_38120),
    .O(net_38172)
  );
  InMux inmux_9_6_38127_38145 (
    .I(net_38127),
    .O(net_38145)
  );
  ClkMux inmux_9_6_5_38192 (
    .I(net_5),
    .O(net_38192)
  );
  SRMux inmux_9_6_9_38193 (
    .I(net_9),
    .O(net_38193)
  );
  InMux inmux_9_7_38236_38269 (
    .I(net_38236),
    .O(net_38269)
  );
  InMux inmux_9_7_38240_38298 (
    .I(net_38240),
    .O(net_38298)
  );
  InMux inmux_9_7_38242_38312 (
    .I(net_38242),
    .O(net_38312)
  );
  InMux inmux_9_7_38244_38280 (
    .I(net_38244),
    .O(net_38280)
  );
  InMux inmux_9_7_38246_38294 (
    .I(net_38246),
    .O(net_38294)
  );
  InMux inmux_9_7_38249_38276 (
    .I(net_38249),
    .O(net_38276)
  );
  InMux inmux_9_7_38253_38304 (
    .I(net_38253),
    .O(net_38304)
  );
  InMux inmux_9_7_38255_38299 (
    .I(net_38255),
    .O(net_38299)
  );
  InMux inmux_9_7_38256_38286 (
    .I(net_38256),
    .O(net_38286)
  );
  ClkMux inmux_9_7_5_38315 (
    .I(net_5),
    .O(net_38315)
  );
  SRMux inmux_9_7_9_38316 (
    .I(net_9),
    .O(net_38316)
  );
  InMux inmux_9_8_38359_38399 (
    .I(net_38359),
    .O(net_38399)
  );
  InMux inmux_9_8_38361_38411 (
    .I(net_38361),
    .O(net_38411)
  );
  InMux inmux_9_8_38363_38423 (
    .I(net_38363),
    .O(net_38423)
  );
  InMux inmux_9_8_38364_38429 (
    .I(net_38364),
    .O(net_38429)
  );
  InMux inmux_9_8_38365_38435 (
    .I(net_38365),
    .O(net_38435)
  );
  InMux inmux_9_8_38368_38404 (
    .I(net_38368),
    .O(net_38404)
  );
  InMux inmux_9_8_38370_38416 (
    .I(net_38370),
    .O(net_38416)
  );
  InMux inmux_9_8_38373_38393 (
    .I(net_38373),
    .O(net_38393)
  );
  InMux inmux_9_8_38375_38392 (
    .I(net_38375),
    .O(net_38392)
  );
  InMux inmux_9_8_38380_38398 (
    .I(net_38380),
    .O(net_38398)
  );
  InMux inmux_9_8_38390_38400 (
    .I(net_38390),
    .O(net_38400)
  );
  InMux inmux_9_8_38396_38406 (
    .I(net_38396),
    .O(net_38406)
  );
  InMux inmux_9_8_38402_38412 (
    .I(net_38402),
    .O(net_38412)
  );
  InMux inmux_9_8_38408_38418 (
    .I(net_38408),
    .O(net_38418)
  );
  InMux inmux_9_8_38414_38424 (
    .I(net_38414),
    .O(net_38424)
  );
  InMux inmux_9_8_38420_38430 (
    .I(net_38420),
    .O(net_38430)
  );
  InMux inmux_9_8_38426_38436 (
    .I(net_38426),
    .O(net_38436)
  );
  ClkMux inmux_9_8_5_38438 (
    .I(net_5),
    .O(net_38438)
  );
  SRMux inmux_9_8_9_38439 (
    .I(net_9),
    .O(net_38439)
  );
  InMux inmux_9_9_38476_38517 (
    .I(net_38476),
    .O(net_38517)
  );
  InMux inmux_9_9_38484_38522 (
    .I(net_38484),
    .O(net_38522)
  );
  InMux inmux_9_9_38485_38559 (
    .I(net_38485),
    .O(net_38559)
  );
  InMux inmux_9_9_38486_38539 (
    .I(net_38486),
    .O(net_38539)
  );
  InMux inmux_9_9_38487_38550 (
    .I(net_38487),
    .O(net_38550)
  );
  InMux inmux_9_9_38491_38532 (
    .I(net_38491),
    .O(net_38532)
  );
  InMux inmux_9_9_38494_38528 (
    .I(net_38494),
    .O(net_38528)
  );
  InMux inmux_9_9_38495_38544 (
    .I(net_38495),
    .O(net_38544)
  );
  ClkMux inmux_9_9_5_38561 (
    .I(net_5),
    .O(net_38561)
  );
  SRMux inmux_9_9_9_38562 (
    .I(net_9),
    .O(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42470_cascademuxed),
    .in3(gnd),
    .lcout(net_38563),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(gnd),
    .in1(net_42475),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38564),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(net_42480),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38565),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(net_42486),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38566),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42500_cascademuxed),
    .in3(gnd),
    .lcout(net_38568),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(gnd),
    .in1(net_42505),
    .in2(net_42506_cascademuxed),
    .in3(gnd),
    .lcout(net_38569),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42515),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42512_cascademuxed),
    .in3(gnd),
    .lcout(net_38570),
    .ltout(),
    .sr(net_42516)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42637),
    .clk(net_42638),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42594),
    .lcout(net_38686),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42637),
    .clk(net_42638),
    .in0(gnd),
    .in1(net_42598),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42637),
    .clk(net_42638),
    .in0(net_42609),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38689),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42615),
    .in1(net_42616),
    .in2(net_42617_cascademuxed),
    .in3(net_42618),
    .lcout(net_38690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42637),
    .clk(net_42638),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42630),
    .lcout(net_38692),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42633),
    .in1(net_42634),
    .in2(net_42635_cascademuxed),
    .in3(net_42636),
    .lcout(net_38693),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42760),
    .clk(net_42761),
    .in0(net_42726),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38811),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42883),
    .clk(net_42884),
    .in0(net_42843),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38933),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42851_cascademuxed),
    .in3(gnd),
    .lcout(net_38934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(net_42961),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39055),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42969),
    .lcout(net_39056),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42980_cascademuxed),
    .in3(gnd),
    .lcout(net_39058),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(net_42985),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39059),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42993),
    .lcout(net_39060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(net_43003),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43129),
    .clk(net_43130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43085_cascademuxed),
    .in3(gnd),
    .lcout(net_39178),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110001000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_43095),
    .in1(net_43096),
    .in2(net_43097_cascademuxed),
    .in3(net_43098),
    .lcout(net_39180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43129),
    .clk(net_43130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43109_cascademuxed),
    .in3(gnd),
    .lcout(net_39182),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43129),
    .clk(net_43130),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_43128),
    .lcout(net_39185),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43252),
    .clk(net_43253),
    .in0(gnd),
    .in1(net_43207),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39301),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43252),
    .clk(net_43253),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_43215),
    .lcout(net_39302),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43252),
    .clk(net_43253),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43226_cascademuxed),
    .in3(gnd),
    .lcout(net_39304),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43252),
    .clk(net_43253),
    .in0(gnd),
    .in1(net_43231),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39305),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43252),
    .clk(net_43253),
    .in0(gnd),
    .in1(net_43237),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39306),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100000111000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_43329),
    .in1(net_43330),
    .in2(net_43331_cascademuxed),
    .in3(net_43332),
    .lcout(net_39424),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43375),
    .clk(net_43376),
    .in0(net_43335),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39425),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_10_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_43341),
    .in1(net_43342),
    .in2(net_43343_cascademuxed),
    .in3(net_43344),
    .lcout(net_39426),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43375),
    .clk(net_43376),
    .in0(net_43353),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39428),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_10_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_43365),
    .in1(net_43366),
    .in2(net_43367_cascademuxed),
    .in3(net_43368),
    .lcout(net_39430),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43375),
    .clk(net_43376),
    .in0(gnd),
    .in1(net_43372),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(net_43452),
    .in1(net_43453),
    .in2(net_43454_cascademuxed),
    .in3(gnd),
    .lcout(net_39547),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100011011000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(net_43458),
    .in1(net_43459),
    .in2(net_43460_cascademuxed),
    .in3(gnd),
    .lcout(net_39548),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43465),
    .in2(net_43466_cascademuxed),
    .in3(net_43467),
    .lcout(net_39549),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111001000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(net_43470),
    .in1(net_43471),
    .in2(gnd),
    .in3(net_43473),
    .lcout(net_39550),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(net_43476),
    .in1(net_43477),
    .in2(net_43478_cascademuxed),
    .in3(gnd),
    .lcout(net_39551),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111111000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43483),
    .in2(net_43484_cascademuxed),
    .in3(net_43485),
    .lcout(net_39552),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(net_43488),
    .in1(net_43489),
    .in2(gnd),
    .in3(net_43491),
    .lcout(net_39553),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43498),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43495),
    .in2(net_43496_cascademuxed),
    .in3(net_43497),
    .lcout(net_39554),
    .ltout(),
    .sr(net_43500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43621),
    .clk(net_43622),
    .in0(net_43581),
    .in1(net_43582),
    .in2(net_43583_cascademuxed),
    .in3(net_43584),
    .lcout(net_39671),
    .ltout(),
    .sr(net_43623)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43621),
    .clk(net_43622),
    .in0(net_43617),
    .in1(net_43618),
    .in2(net_43619_cascademuxed),
    .in3(net_43620),
    .lcout(net_39677),
    .ltout(),
    .sr(net_43623)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_1_0 (
    .carryin(t501),
    .carryout(net_41320),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41322),
    .in2(net_41323_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_1_1 (
    .carryin(net_41320),
    .carryout(net_41326),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41328),
    .in2(net_41329_cascademuxed),
    .in3(net_41330),
    .lcout(net_37416),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_1_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41333),
    .in1(net_41334),
    .in2(gnd),
    .in3(net_41336),
    .lcout(net_37417),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41368),
    .in0(gnd),
    .in1(net_41352),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37420),
    .ltout(),
    .sr(net_41369)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41368),
    .in0(gnd),
    .in1(net_41358),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37421),
    .ltout(),
    .sr(net_41369)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41365_cascademuxed),
    .in3(net_41366),
    .lcout(net_37422),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(net_41485),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37543),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(net_41490),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37544),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(net_41497),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37545),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41504_cascademuxed),
    .in3(gnd),
    .lcout(net_37546),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41511),
    .lcout(net_37547),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41517),
    .lcout(net_37548),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(gnd),
    .in1(net_41521),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37549),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41531),
    .in0(net_41526),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37550),
    .ltout(),
    .sr(net_41532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(net_41608),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37702),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41615_cascademuxed),
    .in3(gnd),
    .lcout(net_37703),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41622),
    .lcout(net_37704),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41627_cascademuxed),
    .in3(gnd),
    .lcout(net_37705),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41633_cascademuxed),
    .in3(gnd),
    .lcout(net_37706),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(net_41637),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37707),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41645_cascademuxed),
    .in3(gnd),
    .lcout(net_37708),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41654),
    .in0(gnd),
    .in1(net_41650),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37709),
    .ltout(),
    .sr(net_41655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41730),
    .in1(net_41731),
    .in2(net_41732_cascademuxed),
    .in3(net_41733),
    .lcout(net_37825),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41776),
    .clk(net_41777),
    .in0(gnd),
    .in1(net_41737),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37826),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41776),
    .clk(net_41777),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41750_cascademuxed),
    .in3(gnd),
    .lcout(net_37828),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41776),
    .clk(net_41777),
    .in0(gnd),
    .in1(net_41761),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41776),
    .clk(net_41777),
    .in0(net_41766),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37831),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_10_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41772),
    .in1(net_41773),
    .in2(net_41774_cascademuxed),
    .in3(net_41775),
    .lcout(net_37832),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41900),
    .in0(net_41859),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37949),
    .ltout(),
    .sr(net_41901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41900),
    .in0(net_41877),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37952),
    .ltout(),
    .sr(net_41901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41900),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41886),
    .lcout(net_37953),
    .ltout(),
    .sr(net_41901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41900),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41892),
    .lcout(net_37954),
    .ltout(),
    .sr(net_41901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_41900),
    .in0(net_41895),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37955),
    .ltout(),
    .sr(net_41901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42022),
    .clk(net_42023),
    .in0(gnd),
    .in1(net_41983),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38072),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42022),
    .clk(net_42023),
    .in0(gnd),
    .in1(net_42001),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38075),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42022),
    .clk(net_42023),
    .in0(net_42018),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38078),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(gnd),
    .in1(net_42100),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38194),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42107_cascademuxed),
    .in3(gnd),
    .lcout(net_38195),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(gnd),
    .in1(net_42118),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38197),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(net_42123),
    .in1(gnd),
    .in2(net_42125_cascademuxed),
    .in3(gnd),
    .lcout(net_38198),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(gnd),
    .in1(net_42130),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38199),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42146),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42144),
    .lcout(net_38201),
    .ltout(),
    .sr(net_42147)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42225),
    .lcout(net_38317),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(net_42229),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38318),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(net_42240),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38320),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42248_cascademuxed),
    .in3(gnd),
    .lcout(net_38321),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42255),
    .lcout(net_38322),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(net_42259),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38323),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_42269),
    .in0(gnd),
    .in1(net_42265),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38324),
    .ltout(),
    .sr(net_42270)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42391),
    .clk(net_42392),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42365_cascademuxed),
    .in3(gnd),
    .lcout(net_38443),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46345),
    .clk(net_46346),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46307_cascademuxed),
    .in3(gnd),
    .lcout(net_42395),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46345),
    .clk(net_46346),
    .in0(gnd),
    .in1(net_46324),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42398),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46345),
    .clk(net_46346),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46343_cascademuxed),
    .in3(gnd),
    .lcout(net_42401),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110001100100),
    .SEQ_MODE(4'b0000)
  ) lc40_11_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46422),
    .in1(net_46423),
    .in2(net_46424_cascademuxed),
    .in3(net_46425),
    .lcout(net_42517),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(net_46429),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42518),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(net_46434),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46437),
    .lcout(net_42519),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46442_cascademuxed),
    .in3(net_46443),
    .lcout(net_42520),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(net_46447),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42521),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46455),
    .lcout(net_42522),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(net_46459),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42523),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46469),
    .in0(gnd),
    .in1(net_46465),
    .in2(gnd),
    .in3(net_46467),
    .lcout(net_42524),
    .ltout(),
    .sr(net_46470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000011001100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(gnd),
    .in1(net_46546),
    .in2(net_46547_cascademuxed),
    .in3(net_46548),
    .lcout(net_42640),
    .ltout(),
    .sr(net_46593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100011011000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(net_46551),
    .in1(net_46552),
    .in2(net_46553_cascademuxed),
    .in3(gnd),
    .lcout(net_42641),
    .ltout(),
    .sr(net_46593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101110001000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(net_46557),
    .in1(net_46558),
    .in2(gnd),
    .in3(net_46560),
    .lcout(net_42642),
    .ltout(),
    .sr(net_46593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101010001010),
    .SEQ_MODE(4'b0000)
  ) lc40_11_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46569),
    .in1(net_46570),
    .in2(net_46571_cascademuxed),
    .in3(net_46572),
    .lcout(net_42644),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(net_46575),
    .in1(net_46576),
    .in2(net_46577_cascademuxed),
    .in3(gnd),
    .lcout(net_42645),
    .ltout(),
    .sr(net_46593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010110000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46680),
    .in1(net_46681),
    .in2(net_46682_cascademuxed),
    .in3(net_46683),
    .lcout(net_42765),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46714),
    .clk(net_46715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46694_cascademuxed),
    .in3(gnd),
    .lcout(net_42767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46794),
    .lcout(net_42886),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46806),
    .lcout(net_42888),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46817_cascademuxed),
    .in3(gnd),
    .lcout(net_42890),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46824),
    .lcout(net_42891),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(net_46834),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42893),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(gnd),
    .in1(net_46915),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43009),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46923),
    .lcout(net_43010),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_11_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46926),
    .in1(net_46927),
    .in2(net_46928_cascademuxed),
    .in3(net_46929),
    .lcout(net_43011),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(net_46938),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43013),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(net_46950),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43015),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110001100100),
    .SEQ_MODE(4'b0000)
  ) lc40_11_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46956),
    .in1(net_46957),
    .in2(net_46958_cascademuxed),
    .in3(net_46959),
    .lcout(net_43016),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47083),
    .clk(net_47084),
    .in0(net_47037),
    .in1(net_47038),
    .in2(net_47039_cascademuxed),
    .in3(gnd),
    .lcout(net_43132),
    .ltout(),
    .sr(net_47085)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110100000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47083),
    .clk(net_47084),
    .in0(net_47043),
    .in1(gnd),
    .in2(net_47045_cascademuxed),
    .in3(net_47046),
    .lcout(net_43133),
    .ltout(),
    .sr(net_47085)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47083),
    .clk(net_47084),
    .in0(net_47055),
    .in1(net_47056),
    .in2(net_47057_cascademuxed),
    .in3(gnd),
    .lcout(net_43135),
    .ltout(),
    .sr(net_47085)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47083),
    .clk(net_47084),
    .in0(gnd),
    .in1(net_47062),
    .in2(net_47063_cascademuxed),
    .in3(net_47064),
    .lcout(net_43136),
    .ltout(),
    .sr(net_47085)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47206),
    .clk(net_47207),
    .in0(gnd),
    .in1(gnd),
    .in2(net_47162_cascademuxed),
    .in3(gnd),
    .lcout(net_43255),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47206),
    .clk(net_47207),
    .in0(gnd),
    .in1(net_47173),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43257),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47206),
    .clk(net_47207),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_47181),
    .lcout(net_43258),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47206),
    .clk(net_47207),
    .in0(gnd),
    .in1(net_47185),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43259),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010001100),
    .SEQ_MODE(4'b0000)
  ) lc40_11_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_47190),
    .in1(net_47191),
    .in2(net_47192_cascademuxed),
    .in3(net_47193),
    .lcout(net_43260),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_11_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_47196),
    .in1(net_47197),
    .in2(net_47198_cascademuxed),
    .in3(net_47199),
    .lcout(net_43261),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47206),
    .clk(net_47207),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_47205),
    .lcout(net_43262),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010010100100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(net_47289),
    .in1(net_47290),
    .in2(net_47291_cascademuxed),
    .in3(net_47292),
    .lcout(net_43379),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110010011000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(net_47295),
    .in1(net_47296),
    .in2(net_47297_cascademuxed),
    .in3(net_47298),
    .lcout(net_43380),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(net_47313),
    .in1(net_47314),
    .in2(net_47315_cascademuxed),
    .in3(net_47316),
    .lcout(net_43383),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101010011000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(net_47325),
    .in1(net_47326),
    .in2(net_47327_cascademuxed),
    .in3(net_47328),
    .lcout(net_43385),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47452),
    .clk(net_47453),
    .in0(gnd),
    .in1(net_47413),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43502),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_1_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45199),
    .in0(gnd),
    .in1(gnd),
    .in2(net_45178_cascademuxed),
    .in3(gnd),
    .lcout(net_41250),
    .ltout(),
    .sr(net_45200)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_2_0 (
    .carryin(t549),
    .carryout(net_45314),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45316),
    .in2(net_45317_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_2_1 (
    .carryin(net_45314),
    .carryout(net_45320),
    .ce(),
    .clk(net_45362),
    .in0(gnd),
    .in1(net_45322),
    .in2(net_45323_cascademuxed),
    .in3(net_45324),
    .lcout(net_41375),
    .ltout(),
    .sr(net_45363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45362),
    .in0(gnd),
    .in1(net_45328),
    .in2(net_45329_cascademuxed),
    .in3(net_45330),
    .lcout(net_41376),
    .ltout(),
    .sr(net_45363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_11_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45340),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41378),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45362),
    .in0(net_45345),
    .in1(gnd),
    .in2(net_45347_cascademuxed),
    .in3(gnd),
    .lcout(net_41379),
    .ltout(),
    .sr(net_45363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45362),
    .in0(gnd),
    .in1(gnd),
    .in2(net_45353_cascademuxed),
    .in3(gnd),
    .lcout(net_41380),
    .ltout(),
    .sr(net_45363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45362),
    .in0(net_45357),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41381),
    .ltout(),
    .sr(net_45363)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_0 (
    .carryin(t552),
    .carryout(net_45437),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45439),
    .in2(net_45440_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_1 (
    .carryin(net_45437),
    .carryout(net_45443),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45445),
    .in2(net_45446_cascademuxed),
    .in3(net_45447),
    .lcout(net_41534),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_2 (
    .carryin(net_45443),
    .carryout(net_45449),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45451),
    .in2(net_45452_cascademuxed),
    .in3(net_45453),
    .lcout(net_41535),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_3 (
    .carryin(net_45449),
    .carryout(net_45455),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45457),
    .in2(net_45458_cascademuxed),
    .in3(net_45459),
    .lcout(net_41536),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_4 (
    .carryin(net_45455),
    .carryout(net_45461),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45463),
    .in2(net_45464_cascademuxed),
    .in3(net_45465),
    .lcout(net_41537),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_5 (
    .carryin(net_45461),
    .carryout(net_45467),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45469),
    .in2(net_45470_cascademuxed),
    .in3(net_45471),
    .lcout(net_41538),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_6 (
    .carryin(net_45467),
    .carryout(net_45473),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45475),
    .in2(net_45476_cascademuxed),
    .in3(net_45477),
    .lcout(net_41539),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_3_7 (
    .carryin(net_45473),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45483),
    .lcout(net_41540),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_4_0 (
    .carryin(t558),
    .carryout(net_45560),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45562),
    .in2(net_45563_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_1 (
    .carryin(net_45560),
    .carryout(net_45566),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45568),
    .in2(net_45569_cascademuxed),
    .in3(net_45570),
    .lcout(net_41657),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_2 (
    .carryin(net_45566),
    .carryout(net_45572),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45574),
    .in2(net_45575_cascademuxed),
    .in3(net_45576),
    .lcout(net_41658),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_3 (
    .carryin(net_45572),
    .carryout(net_45578),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45580),
    .in2(net_45581_cascademuxed),
    .in3(net_45582),
    .lcout(net_41659),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_4 (
    .carryin(net_45578),
    .carryout(net_45584),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45586),
    .in2(net_45587_cascademuxed),
    .in3(net_45588),
    .lcout(net_41660),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_5 (
    .carryin(net_45584),
    .carryout(net_45590),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45592),
    .in2(net_45593_cascademuxed),
    .in3(net_45594),
    .lcout(net_41661),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_6 (
    .carryin(net_45590),
    .carryout(net_45596),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45598),
    .in2(net_45599_cascademuxed),
    .in3(net_45600),
    .lcout(net_41662),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_4_7 (
    .carryin(net_45596),
    .carryout(net_45602),
    .ce(),
    .clk(net_45608),
    .in0(gnd),
    .in1(net_45604),
    .in2(net_45605_cascademuxed),
    .in3(net_45606),
    .lcout(net_41663),
    .ltout(),
    .sr(net_45609)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_0 (
    .carryin(net_45646),
    .carryout(net_45683),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(net_45685),
    .in2(gnd),
    .in3(net_45687),
    .lcout(net_41779),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(gnd),
    .in2(net_45692_cascademuxed),
    .in3(net_45693),
    .lcout(net_41780),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(net_45697),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41781),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(net_45702),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41782),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45711),
    .lcout(net_41783),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(net_45715),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41784),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(net_45720),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41785),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45731),
    .in0(gnd),
    .in1(net_45727),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41786),
    .ltout(),
    .sr(net_45732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45854),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45810),
    .lcout(net_41902),
    .ltout(),
    .sr(net_45855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45854),
    .in0(gnd),
    .in1(net_45814),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41903),
    .ltout(),
    .sr(net_45855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45854),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45834),
    .lcout(net_41906),
    .ltout(),
    .sr(net_45855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_45854),
    .in0(gnd),
    .in1(net_45850),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_41909),
    .ltout(),
    .sr(net_45855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_45976),
    .clk(net_45977),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45933),
    .lcout(net_42025),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_45976),
    .clk(net_45977),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_45957),
    .lcout(net_42029),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_45976),
    .clk(net_45977),
    .in0(net_45960),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42030),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46055_cascademuxed),
    .in3(gnd),
    .lcout(net_42148),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46061_cascademuxed),
    .in3(gnd),
    .lcout(net_42149),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(gnd),
    .in1(net_46066),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42150),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(net_46071),
    .in1(net_46072),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42151),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46079_cascademuxed),
    .in3(gnd),
    .lcout(net_42152),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(gnd),
    .in1(net_46084),
    .in2(gnd),
    .in3(net_46086),
    .lcout(net_42153),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(net_46089),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46092),
    .lcout(net_42154),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46100),
    .in0(net_46095),
    .in1(net_46096),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42155),
    .ltout(),
    .sr(net_46101)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46223),
    .in0(gnd),
    .in1(net_46183),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42272),
    .ltout(),
    .sr(net_46224)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46223),
    .in0(gnd),
    .in1(net_46201),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42275),
    .ltout(),
    .sr(net_46224)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_46223),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46221),
    .lcout(net_42278),
    .ltout(),
    .sr(net_46224)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50177),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50139),
    .lcout(net_46226),
    .ltout(),
    .sr(net_50178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50177),
    .in0(gnd),
    .in1(net_50149),
    .in2(gnd),
    .in3(net_50151),
    .lcout(net_46228),
    .ltout(),
    .sr(net_50178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50177),
    .in0(net_50154),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46229),
    .ltout(),
    .sr(net_50178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50177),
    .in0(net_50166),
    .in1(gnd),
    .in2(net_50168_cascademuxed),
    .in3(gnd),
    .lcout(net_46231),
    .ltout(),
    .sr(net_50178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50177),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50174_cascademuxed),
    .in3(gnd),
    .lcout(net_46232),
    .ltout(),
    .sr(net_50178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(net_50265),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46350),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50274),
    .lcout(net_46351),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50279_cascademuxed),
    .in3(gnd),
    .lcout(net_46352),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50285_cascademuxed),
    .in3(gnd),
    .lcout(net_46353),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50291_cascademuxed),
    .in3(gnd),
    .lcout(net_46354),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50379),
    .lcout(net_46471),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50383),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46472),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101011010000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50394),
    .in1(net_50395),
    .in2(net_50396_cascademuxed),
    .in3(net_50397),
    .lcout(net_46474),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50501_cascademuxed),
    .in3(gnd),
    .lcout(net_46594),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50514),
    .lcout(net_46596),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(net_50517),
    .in1(net_50518),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46597),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(net_50523),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46598),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50532),
    .lcout(net_46599),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50546),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50538),
    .lcout(net_46600),
    .ltout(),
    .sr(net_50547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50622),
    .in1(gnd),
    .in2(net_50624_cascademuxed),
    .in3(net_50625),
    .lcout(net_46717),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100011011000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50628),
    .in1(net_50629),
    .in2(net_50630_cascademuxed),
    .in3(gnd),
    .lcout(net_46718),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111110100000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50640),
    .in1(gnd),
    .in2(net_50642_cascademuxed),
    .in3(net_50643),
    .lcout(net_46720),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(gnd),
    .in1(net_50647),
    .in2(net_50648_cascademuxed),
    .in3(net_50649),
    .lcout(net_46721),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50652),
    .in1(gnd),
    .in2(net_50654_cascademuxed),
    .in3(gnd),
    .lcout(net_46722),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101110001000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50658),
    .in1(net_50659),
    .in2(gnd),
    .in3(net_50661),
    .lcout(net_46723),
    .ltout(),
    .sr(net_50670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50791),
    .clk(net_50792),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50748),
    .lcout(net_46840),
    .ltout(),
    .sr(net_50793)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50751),
    .in1(net_50752),
    .in2(net_50753_cascademuxed),
    .in3(net_50754),
    .lcout(net_46841),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50757),
    .in1(net_50758),
    .in2(net_50759_cascademuxed),
    .in3(net_50760),
    .lcout(net_46842),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50763),
    .in1(net_50764),
    .in2(net_50765_cascademuxed),
    .in3(net_50766),
    .lcout(net_46843),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_50770),
    .in2(net_50771_cascademuxed),
    .in3(net_50772),
    .lcout(net_46844),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50775),
    .in1(net_50776),
    .in2(net_50777_cascademuxed),
    .in3(gnd),
    .lcout(net_46845),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50787),
    .in1(net_50788),
    .in2(net_50789_cascademuxed),
    .in3(net_50790),
    .lcout(net_46847),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50868),
    .in1(net_50869),
    .in2(net_50870_cascademuxed),
    .in3(net_50871),
    .lcout(net_46963),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000011011111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50874),
    .in1(net_50875),
    .in2(net_50876_cascademuxed),
    .in3(net_50877),
    .lcout(net_46964),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50915),
    .in0(net_50880),
    .in1(gnd),
    .in2(net_50882_cascademuxed),
    .in3(gnd),
    .lcout(net_46965),
    .ltout(),
    .sr(net_50916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50915),
    .in0(net_50886),
    .in1(net_50887),
    .in2(net_50888_cascademuxed),
    .in3(net_50889),
    .lcout(net_46966),
    .ltout(),
    .sr(net_50916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_50915),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50894_cascademuxed),
    .in3(gnd),
    .lcout(net_46967),
    .ltout(),
    .sr(net_50916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101010001010),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50898),
    .in1(net_50899),
    .in2(net_50900_cascademuxed),
    .in3(net_50901),
    .lcout(net_46968),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100110010000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50904),
    .in1(net_50905),
    .in2(net_50906_cascademuxed),
    .in3(net_50907),
    .lcout(net_46969),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50910),
    .in1(net_50911),
    .in2(net_50912_cascademuxed),
    .in3(net_50913),
    .lcout(net_46970),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_17_0 (
    .carryin(t636),
    .carryout(t638),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50993_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_1 (
    .carryin(t638),
    .carryout(net_50996),
    .ce(),
    .clk(net_51038),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50999_cascademuxed),
    .in3(net_51000),
    .lcout(net_47087),
    .ltout(),
    .sr(net_51039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_51038),
    .in0(net_51003),
    .in1(gnd),
    .in2(gnd),
    .in3(net_51006),
    .lcout(net_47088),
    .ltout(),
    .sr(net_51039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_51038),
    .in0(gnd),
    .in1(gnd),
    .in2(net_51011_cascademuxed),
    .in3(gnd),
    .lcout(net_47089),
    .ltout(),
    .sr(net_51039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_12_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_51016),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47090),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_51038),
    .in0(net_51027),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47092),
    .ltout(),
    .sr(net_51039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_51038),
    .in0(gnd),
    .in1(gnd),
    .in2(net_51035_cascademuxed),
    .in3(gnd),
    .lcout(net_47093),
    .ltout(),
    .sr(net_51039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51160),
    .clk(net_51161),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_51129),
    .lcout(net_47211),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51160),
    .clk(net_51161),
    .in0(gnd),
    .in1(net_51139),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47213),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51283),
    .clk(net_51284),
    .in0(net_51255),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47335),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_1_0 (
    .carryin(t591),
    .carryout(t593),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_48985_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0001000101000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_1_1 (
    .carryin(t593),
    .carryout(net_48988),
    .ce(net_49029),
    .clk(net_49030),
    .in0(net_48989),
    .in1(net_48990),
    .in2(gnd),
    .in3(net_48992),
    .lcout(net_45078),
    .ltout(),
    .sr(net_49031)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000010101010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_1_2 (
    .carryin(net_48988),
    .carryout(net_48994),
    .ce(net_49029),
    .clk(net_49030),
    .in0(net_48995),
    .in1(gnd),
    .in2(net_48997_cascademuxed),
    .in3(net_48998),
    .lcout(net_45079),
    .ltout(),
    .sr(net_49031)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0001000101000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_1_3 (
    .carryin(net_48994),
    .carryout(net_49000),
    .ce(net_49029),
    .clk(net_49030),
    .in0(net_49001),
    .in1(net_49002),
    .in2(gnd),
    .in3(net_49004),
    .lcout(net_45080),
    .ltout(),
    .sr(net_49031)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100110000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_1_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49029),
    .clk(net_49030),
    .in0(gnd),
    .in1(net_49008),
    .in2(net_49009_cascademuxed),
    .in3(net_49010),
    .lcout(net_45081),
    .ltout(),
    .sr(net_49031)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49148_cascademuxed),
    .in3(gnd),
    .lcout(net_45205),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49193),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49155),
    .lcout(net_45206),
    .ltout(),
    .sr(net_49194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_12_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49158),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45207),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49193),
    .in0(net_49164),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45208),
    .ltout(),
    .sr(net_49194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49193),
    .in0(net_49170),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45209),
    .ltout(),
    .sr(net_49194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49193),
    .in0(gnd),
    .in1(net_49183),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45211),
    .ltout(),
    .sr(net_49194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_3_0 (
    .carryin(t650),
    .carryout(t653),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49271_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_3_1 (
    .carryin(t653),
    .carryout(t654),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_49276),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_3_2 (
    .carryin(t654),
    .carryout(t655),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_49282),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_3_3 (
    .carryin(t655),
    .carryout(net_49286),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49289_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011110011),
    .SEQ_MODE(4'b0000)
  ) lc40_12_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_49294),
    .in2(net_49295_cascademuxed),
    .in3(net_49296),
    .lcout(net_45368),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49316),
    .in0(net_49299),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45369),
    .ltout(),
    .sr(net_49317)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49316),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49308),
    .lcout(net_45370),
    .ltout(),
    .sr(net_49317)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49316),
    .in0(gnd),
    .in1(net_49312),
    .in2(gnd),
    .in3(net_49314),
    .lcout(net_45371),
    .ltout(),
    .sr(net_49317)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49438),
    .clk(net_49439),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49395),
    .lcout(net_45487),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_12_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49398),
    .in1(net_49399),
    .in2(net_49400_cascademuxed),
    .in3(net_49401),
    .lcout(net_45488),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49438),
    .clk(net_49439),
    .in0(gnd),
    .in1(net_49405),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45489),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_12_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49410),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45490),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49438),
    .clk(net_49439),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49418_cascademuxed),
    .in3(gnd),
    .lcout(net_45491),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49422),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49425),
    .lcout(net_45492),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010110000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49428),
    .in1(net_49429),
    .in2(net_49430_cascademuxed),
    .in3(net_49431),
    .lcout(net_45493),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_49435),
    .in2(gnd),
    .in3(net_49437),
    .lcout(net_45494),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49561),
    .clk(net_49562),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49517_cascademuxed),
    .in3(gnd),
    .lcout(net_45610),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49561),
    .clk(net_49562),
    .in0(net_49527),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45612),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49561),
    .clk(net_49562),
    .in0(gnd),
    .in1(net_49546),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45615),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49561),
    .clk(net_49562),
    .in0(gnd),
    .in1(net_49552),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45616),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49640_cascademuxed),
    .in3(gnd),
    .lcout(net_45733),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(net_49645),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45734),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49653),
    .lcout(net_45735),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(net_49656),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45736),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(net_49663),
    .in2(gnd),
    .in3(net_49665),
    .lcout(net_45737),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49670_cascademuxed),
    .in3(net_49671),
    .lcout(net_45738),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(net_49674),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49677),
    .lcout(net_45739),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_49685),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_49683),
    .lcout(net_45740),
    .ltout(),
    .sr(net_49686)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49807),
    .clk(net_49808),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49763_cascademuxed),
    .in3(gnd),
    .lcout(net_45856),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49807),
    .clk(net_49808),
    .in0(net_49767),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45857),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_12_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49779),
    .in1(net_49780),
    .in2(net_49781_cascademuxed),
    .in3(net_49782),
    .lcout(net_45859),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49807),
    .clk(net_49808),
    .in0(net_49785),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45860),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49807),
    .clk(net_49808),
    .in0(net_49797),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45862),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49807),
    .clk(net_49808),
    .in0(gnd),
    .in1(net_49804),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45863),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49930),
    .clk(net_49931),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49886_cascademuxed),
    .in3(gnd),
    .lcout(net_45979),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49930),
    .clk(net_49931),
    .in0(gnd),
    .in1(net_49909),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45983),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49930),
    .clk(net_49931),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49916_cascademuxed),
    .in3(gnd),
    .lcout(net_45984),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49930),
    .clk(net_49931),
    .in0(gnd),
    .in1(net_49927),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45986),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50053),
    .clk(net_50054),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50010),
    .lcout(net_46102),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50053),
    .clk(net_50054),
    .in0(gnd),
    .in1(net_50038),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46107),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50053),
    .clk(net_50054),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50046),
    .lcout(net_46108),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53961),
    .in1(net_53962),
    .in2(net_53963_cascademuxed),
    .in3(net_53964),
    .lcout(net_50056),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54007),
    .clk(net_54008),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53969_cascademuxed),
    .in3(gnd),
    .lcout(net_50057),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54007),
    .clk(net_54008),
    .in0(gnd),
    .in1(net_53974),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50058),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_13_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53985),
    .in1(net_53986),
    .in2(net_53987_cascademuxed),
    .in3(net_53988),
    .lcout(net_50060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54007),
    .clk(net_54008),
    .in0(net_53991),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50061),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54130),
    .clk(net_54131),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54093),
    .lcout(net_50180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54130),
    .clk(net_54131),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54099),
    .lcout(net_50181),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54108),
    .in1(net_54109),
    .in2(net_54110_cascademuxed),
    .in3(net_54111),
    .lcout(net_50183),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54130),
    .clk(net_54131),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54116_cascademuxed),
    .in3(gnd),
    .lcout(net_50184),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54130),
    .clk(net_54131),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54122_cascademuxed),
    .in3(gnd),
    .lcout(net_50185),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(net_54207),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50302),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54216),
    .lcout(net_50303),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(net_54220),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50304),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54228),
    .lcout(net_50305),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(net_54232),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50306),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54240),
    .lcout(net_50307),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54245_cascademuxed),
    .in3(gnd),
    .lcout(net_50308),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54251_cascademuxed),
    .in3(gnd),
    .lcout(net_50309),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(net_54331),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50425),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011011000100),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54336),
    .in1(net_54337),
    .in2(net_54338_cascademuxed),
    .in3(net_54339),
    .lcout(net_50426),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54345),
    .lcout(net_50427),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54351),
    .lcout(net_50428),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54354),
    .in1(net_54355),
    .in2(net_54356_cascademuxed),
    .in3(net_54357),
    .lcout(net_50429),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(net_54360),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50430),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54366),
    .in1(net_54367),
    .in2(net_54368_cascademuxed),
    .in3(net_54369),
    .lcout(net_50431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54372),
    .in1(net_54373),
    .in2(net_54374_cascademuxed),
    .in3(net_54375),
    .lcout(net_50432),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(net_54453),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54459),
    .in1(gnd),
    .in2(net_54461_cascademuxed),
    .in3(gnd),
    .lcout(net_50549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111011101110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54465),
    .in1(net_54466),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(net_54471),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50551),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(gnd),
    .in1(net_54478),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50552),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54486),
    .lcout(net_50553),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54491_cascademuxed),
    .in3(gnd),
    .lcout(net_50554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101011010000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54495),
    .in1(net_54496),
    .in2(net_54497_cascademuxed),
    .in3(net_54498),
    .lcout(net_50555),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101011111010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54576),
    .in1(gnd),
    .in2(net_54578_cascademuxed),
    .in3(gnd),
    .lcout(net_50671),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54582),
    .in1(gnd),
    .in2(net_54584_cascademuxed),
    .in3(net_54585),
    .lcout(net_50672),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54588),
    .in1(net_54589),
    .in2(net_54590_cascademuxed),
    .in3(net_54591),
    .lcout(net_50673),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54603),
    .lcout(net_50675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(gnd),
    .in1(net_54607),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50676),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54615),
    .lcout(net_50677),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54620_cascademuxed),
    .in3(gnd),
    .lcout(net_50678),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_16_0 (
    .carryin(t686),
    .carryout(t688),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_54700),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_1 (
    .carryin(t688),
    .carryout(net_54704),
    .ce(),
    .clk(net_54746),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54707_cascademuxed),
    .in3(net_54708),
    .lcout(net_50795),
    .ltout(),
    .sr(net_54747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_54746),
    .in0(net_54711),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54714),
    .lcout(net_50796),
    .ltout(),
    .sr(net_54747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54719_cascademuxed),
    .in3(net_54720),
    .lcout(net_50797),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_54746),
    .in0(net_54723),
    .in1(net_54724),
    .in2(net_54725_cascademuxed),
    .in3(net_54726),
    .lcout(net_50798),
    .ltout(),
    .sr(net_54747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100101011001010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54729),
    .in1(net_54730),
    .in2(net_54731_cascademuxed),
    .in3(gnd),
    .lcout(net_50799),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000100001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54735),
    .in1(net_54736),
    .in2(net_54737_cascademuxed),
    .in3(net_54738),
    .lcout(net_50800),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54742),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50801),
    .ltout(),
    .sr(net_54747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_13_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54828),
    .in1(net_54829),
    .in2(gnd),
    .in3(net_54831),
    .lcout(net_50918),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54842_cascademuxed),
    .in3(gnd),
    .lcout(net_50920),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54847),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50921),
    .ltout(),
    .sr(net_54870)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000100001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54852),
    .in1(net_54853),
    .in2(net_54854_cascademuxed),
    .in3(net_54855),
    .lcout(net_50922),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54865),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50924),
    .ltout(),
    .sr(net_54870)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54945),
    .in1(net_54946),
    .in2(net_54947_cascademuxed),
    .in3(net_54948),
    .lcout(net_51040),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54951),
    .in1(net_54952),
    .in2(net_54953_cascademuxed),
    .in3(net_54954),
    .lcout(net_51041),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010111100000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54957),
    .in1(net_54958),
    .in2(net_54959_cascademuxed),
    .in3(net_54960),
    .lcout(net_51042),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54963),
    .in1(net_54964),
    .in2(net_54965_cascademuxed),
    .in3(net_54966),
    .lcout(net_51043),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54975),
    .in1(net_54976),
    .in2(net_54977_cascademuxed),
    .in3(net_54978),
    .lcout(net_51045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54981),
    .in1(net_54982),
    .in2(net_54983_cascademuxed),
    .in3(net_54984),
    .lcout(net_51046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(net_54987),
    .in1(net_54988),
    .in2(net_54989_cascademuxed),
    .in3(net_54990),
    .lcout(net_51047),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55114),
    .clk(net_55115),
    .in0(net_55110),
    .in1(net_55111),
    .in2(net_55112_cascademuxed),
    .in3(net_55113),
    .lcout(net_51170),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_52861),
    .in0(net_52832),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_48911),
    .ltout(),
    .sr(net_52862)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_52846_cascademuxed),
    .in3(net_52847),
    .lcout(net_48913),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_52850),
    .in1(net_52851),
    .in2(net_52852_cascademuxed),
    .in3(gnd),
    .lcout(net_48914),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_52977),
    .in1(gnd),
    .in2(gnd),
    .in3(net_52980),
    .lcout(net_49036),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_52984),
    .in2(net_52985_cascademuxed),
    .in3(net_52986),
    .lcout(net_49037),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53023),
    .clk(net_53024),
    .in0(gnd),
    .in1(net_52990),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49038),
    .ltout(),
    .sr(net_53025)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001010101),
    .SEQ_MODE(4'b0000)
  ) lc40_13_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_52995),
    .in1(gnd),
    .in2(gnd),
    .in3(net_52998),
    .lcout(net_49039),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53023),
    .clk(net_53024),
    .in0(gnd),
    .in1(net_53002),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49040),
    .ltout(),
    .sr(net_53025)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(gnd),
    .in1(net_53101),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49195),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53109),
    .lcout(net_49196),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(net_53112),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49197),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53126_cascademuxed),
    .in3(net_53127),
    .lcout(net_49199),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(gnd),
    .in1(net_53131),
    .in2(net_53132_cascademuxed),
    .in3(gnd),
    .lcout(net_49200),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53147),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53138_cascademuxed),
    .in3(gnd),
    .lcout(net_49201),
    .ltout(),
    .sr(net_53148)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53142),
    .in1(gnd),
    .in2(net_53144_cascademuxed),
    .in3(net_53145),
    .lcout(net_49202),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(net_53223),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49318),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53231_cascademuxed),
    .in3(gnd),
    .lcout(net_49319),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(net_53235),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49320),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53241),
    .in1(net_53242),
    .in2(gnd),
    .in3(net_53244),
    .lcout(net_49321),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(gnd),
    .in1(net_53248),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49322),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53256),
    .lcout(net_49323),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53259),
    .in1(net_53260),
    .in2(net_53261_cascademuxed),
    .in3(net_53262),
    .lcout(net_49324),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_53270),
    .in0(net_53265),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53268),
    .lcout(net_49325),
    .ltout(),
    .sr(net_53271)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53392),
    .clk(net_53393),
    .in0(net_53346),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49441),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53392),
    .clk(net_53393),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53354_cascademuxed),
    .in3(gnd),
    .lcout(net_49442),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53392),
    .clk(net_53393),
    .in0(gnd),
    .in1(net_53377),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49446),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53392),
    .clk(net_53393),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53384_cascademuxed),
    .in3(gnd),
    .lcout(net_49447),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53472),
    .lcout(net_49564),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(net_53475),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49565),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53484),
    .lcout(net_49566),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(net_53487),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49567),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010001100),
    .SEQ_MODE(4'b0000)
  ) lc40_13_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53493),
    .in1(net_53494),
    .in2(net_53495_cascademuxed),
    .in3(net_53496),
    .lcout(net_49568),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(gnd),
    .in1(net_53500),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49569),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(net_53505),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49570),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53515),
    .clk(net_53516),
    .in0(gnd),
    .in1(net_53512),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49571),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53595),
    .lcout(net_49687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53600_cascademuxed),
    .in3(gnd),
    .lcout(net_49688),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53604),
    .in1(net_53605),
    .in2(net_53606_cascademuxed),
    .in3(net_53607),
    .lcout(net_49689),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(net_53610),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(net_53616),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49691),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53624_cascademuxed),
    .in3(gnd),
    .lcout(net_49692),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53638),
    .clk(net_53639),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53630_cascademuxed),
    .in3(gnd),
    .lcout(net_49693),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001110001000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53634),
    .in1(net_53635),
    .in2(net_53636_cascademuxed),
    .in3(net_53637),
    .lcout(net_49694),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53715),
    .in1(net_53716),
    .in2(net_53717_cascademuxed),
    .in3(net_53718),
    .lcout(net_49810),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101010001010),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53721),
    .in1(net_53722),
    .in2(net_53723_cascademuxed),
    .in3(net_53724),
    .lcout(net_49811),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53761),
    .clk(net_53762),
    .in0(net_53727),
    .in1(net_53728),
    .in2(net_53729_cascademuxed),
    .in3(gnd),
    .lcout(net_49812),
    .ltout(),
    .sr(net_53763)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111110100000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53761),
    .clk(net_53762),
    .in0(net_53739),
    .in1(gnd),
    .in2(net_53741_cascademuxed),
    .in3(net_53742),
    .lcout(net_49814),
    .ltout(),
    .sr(net_53763)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53761),
    .clk(net_53762),
    .in0(net_53745),
    .in1(net_53746),
    .in2(net_53747_cascademuxed),
    .in3(gnd),
    .lcout(net_49815),
    .ltout(),
    .sr(net_53763)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53761),
    .clk(net_53762),
    .in0(net_53751),
    .in1(gnd),
    .in2(net_53753_cascademuxed),
    .in3(net_53754),
    .lcout(net_49816),
    .ltout(),
    .sr(net_53763)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101110001000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53761),
    .clk(net_53762),
    .in0(net_53757),
    .in1(net_53758),
    .in2(gnd),
    .in3(net_53760),
    .lcout(net_49817),
    .ltout(),
    .sr(net_53763)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53852_cascademuxed),
    .in3(gnd),
    .lcout(net_49935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53871),
    .lcout(net_49938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(gnd),
    .in1(net_57792),
    .in2(gnd),
    .in3(net_57794),
    .lcout(net_53887),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(net_57797),
    .in1(gnd),
    .in2(net_57799_cascademuxed),
    .in3(gnd),
    .lcout(net_53888),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(net_57803),
    .in1(net_57804),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53889),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(net_57809),
    .in1(net_57810),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53890),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57817_cascademuxed),
    .in3(gnd),
    .lcout(net_53891),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(net_57821),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57824),
    .lcout(net_53892),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(gnd),
    .in1(net_57828),
    .in2(gnd),
    .in3(net_57830),
    .lcout(net_53893),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57838),
    .in0(gnd),
    .in1(net_57834),
    .in2(net_57835_cascademuxed),
    .in3(gnd),
    .lcout(net_53894),
    .ltout(),
    .sr(net_57839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(net_57914),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54010),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57934_cascademuxed),
    .in3(gnd),
    .lcout(net_54013),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(gnd),
    .in1(net_57939),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54014),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57959),
    .lcout(net_54017),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58084),
    .in0(gnd),
    .in1(net_58062),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54137),
    .ltout(),
    .sr(net_58085)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(net_58160),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54256),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(gnd),
    .in1(net_58167),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54257),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58174_cascademuxed),
    .in3(gnd),
    .lcout(net_54258),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111010101110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(net_58178),
    .in1(net_58179),
    .in2(net_58180_cascademuxed),
    .in3(gnd),
    .lcout(net_54259),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58186_cascademuxed),
    .in3(gnd),
    .lcout(net_54260),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58193),
    .lcout(net_54261),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100100011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(net_58196),
    .in1(net_58197),
    .in2(net_58198_cascademuxed),
    .in3(net_58199),
    .lcout(net_54262),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58207),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58204_cascademuxed),
    .in3(gnd),
    .lcout(net_54263),
    .ltout(),
    .sr(net_58208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(gnd),
    .in1(net_58284),
    .in2(net_58285_cascademuxed),
    .in3(gnd),
    .lcout(net_54379),
    .ltout(),
    .sr(net_58331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(gnd),
    .in1(net_58296),
    .in2(gnd),
    .in3(net_58298),
    .lcout(net_54381),
    .ltout(),
    .sr(net_58331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(net_58307),
    .in1(net_58308),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54383),
    .ltout(),
    .sr(net_58331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(net_58313),
    .in1(net_58314),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54384),
    .ltout(),
    .sr(net_58331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58319),
    .in1(net_58320),
    .in2(net_58321_cascademuxed),
    .in3(net_58322),
    .lcout(net_54385),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(net_58325),
    .in1(gnd),
    .in2(net_58327_cascademuxed),
    .in3(gnd),
    .lcout(net_54386),
    .ltout(),
    .sr(net_58331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58407),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54502),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111101110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58412),
    .in1(net_58413),
    .in2(gnd),
    .in3(net_58415),
    .lcout(net_54503),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58453),
    .in0(gnd),
    .in1(net_58419),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54504),
    .ltout(),
    .sr(net_58454)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58427),
    .lcout(net_54505),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58453),
    .in0(gnd),
    .in1(net_58431),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54506),
    .ltout(),
    .sr(net_58454)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58436),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54507),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58444_cascademuxed),
    .in3(gnd),
    .lcout(net_54508),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58449),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54509),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_0 (
    .carryin(t744),
    .carryout(t746),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58531_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_1 (
    .carryin(t746),
    .carryout(net_58534),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58536),
    .in2(net_58537_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_2 (
    .carryin(net_58534),
    .carryout(net_58540),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58542),
    .in2(net_58543_cascademuxed),
    .in3(net_58544),
    .lcout(net_54627),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_3 (
    .carryin(net_58540),
    .carryout(net_58546),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58548),
    .in2(net_58549_cascademuxed),
    .in3(net_58550),
    .lcout(net_54628),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_4 (
    .carryin(net_58546),
    .carryout(net_58552),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58554),
    .in2(net_58555_cascademuxed),
    .in3(net_58556),
    .lcout(net_54629),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_5 (
    .carryin(net_58552),
    .carryout(net_58558),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58560),
    .in2(net_58561_cascademuxed),
    .in3(net_58562),
    .lcout(net_54630),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_6 (
    .carryin(net_58558),
    .carryout(net_58564),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58566),
    .in2(net_58567_cascademuxed),
    .in3(net_58568),
    .lcout(net_54631),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_7 (
    .carryin(net_58564),
    .carryout(net_58570),
    .ce(),
    .clk(net_58576),
    .in0(gnd),
    .in1(net_58572),
    .in2(net_58573_cascademuxed),
    .in3(net_58574),
    .lcout(net_54632),
    .ltout(),
    .sr(net_58577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_14_17_0 (
    .carryin(net_58614),
    .carryout(net_58651),
    .ce(),
    .clk(net_58699),
    .in0(gnd),
    .in1(net_58653),
    .in2(net_58654_cascademuxed),
    .in3(net_58655),
    .lcout(net_54748),
    .ltout(),
    .sr(net_58700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b1000)
  ) lc40_14_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58699),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58661),
    .lcout(net_54749),
    .ltout(),
    .sr(net_58700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58665),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54750),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58672_cascademuxed),
    .in3(gnd),
    .lcout(net_54751),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58699),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58685),
    .lcout(net_54753),
    .ltout(),
    .sr(net_58700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_58699),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58690_cascademuxed),
    .in3(gnd),
    .lcout(net_54754),
    .ltout(),
    .sr(net_58700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58697),
    .lcout(net_54755),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58775),
    .in1(net_58776),
    .in2(net_58777_cascademuxed),
    .in3(gnd),
    .lcout(net_54871),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58781),
    .in1(net_58782),
    .in2(net_58783_cascademuxed),
    .in3(gnd),
    .lcout(net_54872),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000101010000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58787),
    .in1(net_58788),
    .in2(net_58789_cascademuxed),
    .in3(net_58790),
    .lcout(net_54873),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000011001100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(gnd),
    .in1(net_58794),
    .in2(net_58795_cascademuxed),
    .in3(net_58796),
    .lcout(net_54874),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(gnd),
    .in1(net_58806),
    .in2(net_58807_cascademuxed),
    .in3(net_58808),
    .lcout(net_54876),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100010010000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58811),
    .in1(net_58812),
    .in2(net_58813_cascademuxed),
    .in3(net_58814),
    .lcout(net_54877),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58817),
    .in1(net_58818),
    .in2(net_58819_cascademuxed),
    .in3(net_58820),
    .lcout(net_54878),
    .ltout(),
    .sr(net_58823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110011101100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58944),
    .clk(net_58945),
    .in0(net_58916),
    .in1(net_58917),
    .in2(net_58918_cascademuxed),
    .in3(net_58919),
    .lcout(net_54997),
    .ltout(),
    .sr(net_58946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_56682_cascademuxed),
    .in3(net_56683),
    .lcout(net_52745),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56853),
    .clk(net_56854),
    .in0(gnd),
    .in1(gnd),
    .in2(net_56809_cascademuxed),
    .in3(gnd),
    .lcout(net_52867),
    .ltout(),
    .sr(net_56855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56853),
    .clk(net_56854),
    .in0(gnd),
    .in1(net_56820),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_52869),
    .ltout(),
    .sr(net_56855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_56826),
    .in2(net_56827_cascademuxed),
    .in3(net_56828),
    .lcout(net_52870),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56853),
    .clk(net_56854),
    .in0(gnd),
    .in1(gnd),
    .in2(net_56845_cascademuxed),
    .in3(gnd),
    .lcout(net_52873),
    .ltout(),
    .sr(net_56855)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56976),
    .clk(net_56977),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_56969),
    .lcout(net_53032),
    .ltout(),
    .sr(net_56978)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56976),
    .clk(net_56977),
    .in0(net_56972),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53033),
    .ltout(),
    .sr(net_56978)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57055_cascademuxed),
    .in3(gnd),
    .lcout(net_53149),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57065),
    .in1(net_57066),
    .in2(net_57067_cascademuxed),
    .in3(gnd),
    .lcout(net_53151),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(net_57071),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53152),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57079_cascademuxed),
    .in3(gnd),
    .lcout(net_53153),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(net_57083),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53154),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(net_57089),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53155),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(gnd),
    .in1(net_57096),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53156),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_14_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57176),
    .in1(net_57177),
    .in2(net_57178_cascademuxed),
    .in3(net_57179),
    .lcout(net_53272),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57222),
    .clk(net_57223),
    .in0(gnd),
    .in1(net_57183),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53273),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57222),
    .clk(net_57223),
    .in0(net_57188),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53274),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57222),
    .clk(net_57223),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57197),
    .lcout(net_53275),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100101011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57200),
    .in1(net_57201),
    .in2(net_57202_cascademuxed),
    .in3(net_57203),
    .lcout(net_53276),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57206),
    .in1(net_57207),
    .in2(net_57208_cascademuxed),
    .in3(net_57209),
    .lcout(net_53277),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57222),
    .clk(net_57223),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57214_cascademuxed),
    .in3(gnd),
    .lcout(net_53278),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57222),
    .clk(net_57223),
    .in0(net_57218),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53279),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57346),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57302),
    .lcout(net_53395),
    .ltout(),
    .sr(net_57347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57305),
    .in1(net_57306),
    .in2(net_57307_cascademuxed),
    .in3(net_57308),
    .lcout(net_53396),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_14_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57317),
    .in1(net_57318),
    .in2(net_57319_cascademuxed),
    .in3(net_57320),
    .lcout(net_53398),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57346),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57325_cascademuxed),
    .in3(net_57326),
    .lcout(net_53399),
    .ltout(),
    .sr(net_57347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57346),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57332),
    .lcout(net_53400),
    .ltout(),
    .sr(net_57347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57346),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57337_cascademuxed),
    .in3(gnd),
    .lcout(net_53401),
    .ltout(),
    .sr(net_57347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010001100),
    .SEQ_MODE(4'b0000)
  ) lc40_14_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57341),
    .in1(net_57342),
    .in2(net_57343_cascademuxed),
    .in3(net_57344),
    .lcout(net_53402),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57469),
    .in0(gnd),
    .in1(net_57429),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53519),
    .ltout(),
    .sr(net_57470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57469),
    .in0(net_57440),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53521),
    .ltout(),
    .sr(net_57470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57469),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57455),
    .lcout(net_53523),
    .ltout(),
    .sr(net_57470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57460_cascademuxed),
    .in3(gnd),
    .lcout(net_53524),
    .ltout(),
    .sr(net_57470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57469),
    .in0(gnd),
    .in1(net_57465),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53525),
    .ltout(),
    .sr(net_57470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57547_cascademuxed),
    .in3(gnd),
    .lcout(net_53641),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(gnd),
    .in1(net_57552),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53642),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57559_cascademuxed),
    .in3(gnd),
    .lcout(net_53643),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(net_57563),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53644),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(gnd),
    .in1(net_57570),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53645),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(gnd),
    .in1(net_57576),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53646),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57581),
    .in1(net_57582),
    .in2(net_57583_cascademuxed),
    .in3(net_57584),
    .lcout(net_53647),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_57592),
    .in0(net_57587),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53648),
    .ltout(),
    .sr(net_57593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57714),
    .clk(net_57715),
    .in0(net_57668),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53764),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57714),
    .clk(net_57715),
    .in0(gnd),
    .in1(net_57675),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53765),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57704),
    .in1(net_57705),
    .in2(net_57706_cascademuxed),
    .in3(net_57707),
    .lcout(net_53770),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_0 (
    .carryin(t784),
    .carryout(t786),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61622),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0001000101000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_10_1 (
    .carryin(t786),
    .carryout(net_61626),
    .ce(net_61667),
    .clk(net_61668),
    .in0(net_61627),
    .in1(net_61628),
    .in2(gnd),
    .in3(net_61630),
    .lcout(net_57718),
    .ltout(),
    .sr(net_61669)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0001000101000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_10_2 (
    .carryin(net_61626),
    .carryout(net_61632),
    .ce(net_61667),
    .clk(net_61668),
    .in0(net_61633),
    .in1(net_61634),
    .in2(gnd),
    .in3(net_61636),
    .lcout(net_57719),
    .ltout(),
    .sr(net_61669)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100001010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61667),
    .clk(net_61668),
    .in0(net_61639),
    .in1(gnd),
    .in2(net_61641_cascademuxed),
    .in3(net_61642),
    .lcout(net_57720),
    .ltout(),
    .sr(net_61669)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b1000)
  ) lc40_15_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61667),
    .clk(net_61668),
    .in0(net_61657),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57723),
    .ltout(),
    .sr(net_61669)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111001100),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61664),
    .in2(gnd),
    .in3(net_61666),
    .lcout(net_57724),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61744),
    .in1(gnd),
    .in2(net_61746_cascademuxed),
    .in3(net_61747),
    .lcout(net_57840),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61751),
    .in2(net_61752_cascademuxed),
    .in3(net_61753),
    .lcout(net_57841),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(net_61756),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57842),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61765),
    .lcout(net_57843),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61769),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57844),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61776_cascademuxed),
    .in3(gnd),
    .lcout(net_57845),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(net_61780),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57846),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61791),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61788_cascademuxed),
    .in3(gnd),
    .lcout(net_57847),
    .ltout(),
    .sr(net_61792)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61869_cascademuxed),
    .in3(net_61870),
    .lcout(net_57963),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61874),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57964),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61882),
    .lcout(net_57965),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61887_cascademuxed),
    .in3(gnd),
    .lcout(net_57966),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(net_61891),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57967),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61899_cascademuxed),
    .in3(gnd),
    .lcout(net_57968),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(net_61903),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57969),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61910),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57970),
    .ltout(),
    .sr(net_61915)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_0 (
    .carryin(t791),
    .carryout(net_61989),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61991),
    .in2(net_61992_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_1 (
    .carryin(net_61989),
    .carryout(net_61995),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(net_61997),
    .in2(gnd),
    .in3(net_61999),
    .lcout(net_58087),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_2 (
    .carryin(net_61995),
    .carryout(net_62001),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62004_cascademuxed),
    .in3(net_62005),
    .lcout(net_58088),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_3 (
    .carryin(net_62001),
    .carryout(net_62007),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62010_cascademuxed),
    .in3(net_62011),
    .lcout(net_58089),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_4 (
    .carryin(net_62007),
    .carryout(net_62013),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(net_62015),
    .in2(gnd),
    .in3(net_62017),
    .lcout(net_58090),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_5 (
    .carryin(net_62013),
    .carryout(net_62019),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(net_62021),
    .in2(gnd),
    .in3(net_62023),
    .lcout(net_58091),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_13_6 (
    .carryin(net_62019),
    .carryout(net_62025),
    .ce(),
    .clk(net_62037),
    .in0(gnd),
    .in1(net_62027),
    .in2(gnd),
    .in3(net_62029),
    .lcout(net_58092),
    .ltout(),
    .sr(net_62038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_7 (
    .carryin(net_62025),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62035),
    .lcout(net_58093),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62115_cascademuxed),
    .in3(gnd),
    .lcout(net_58209),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(net_62119),
    .in1(gnd),
    .in2(net_62121_cascademuxed),
    .in3(gnd),
    .lcout(net_58210),
    .ltout(),
    .sr(net_62161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62127_cascademuxed),
    .in3(net_62128),
    .lcout(net_58211),
    .ltout(),
    .sr(net_62161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(net_62131),
    .in1(gnd),
    .in2(net_62133_cascademuxed),
    .in3(gnd),
    .lcout(net_58212),
    .ltout(),
    .sr(net_62161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(gnd),
    .in1(net_62138),
    .in2(gnd),
    .in3(net_62140),
    .lcout(net_58213),
    .ltout(),
    .sr(net_62161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62144),
    .in2(net_62145_cascademuxed),
    .in3(gnd),
    .lcout(net_58214),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(gnd),
    .in1(net_62150),
    .in2(gnd),
    .in3(net_62152),
    .lcout(net_58215),
    .ltout(),
    .sr(net_62161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111001100),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62156),
    .in2(gnd),
    .in3(net_62158),
    .lcout(net_58216),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(net_62236),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58332),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62245),
    .lcout(net_58333),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62250_cascademuxed),
    .in3(gnd),
    .lcout(net_58334),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62256_cascademuxed),
    .in3(gnd),
    .lcout(net_58335),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(gnd),
    .in1(net_62261),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58336),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(net_62272),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58338),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62283),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62280_cascademuxed),
    .in3(gnd),
    .lcout(net_58339),
    .ltout(),
    .sr(net_62284)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_0 (
    .carryin(t802),
    .carryout(t804),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62361_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_1 (
    .carryin(t804),
    .carryout(net_62364),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62366),
    .in2(net_62367_cascademuxed),
    .in3(net_62368),
    .lcout(net_58456),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_2 (
    .carryin(net_62364),
    .carryout(net_62370),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62372),
    .in2(net_62373_cascademuxed),
    .in3(net_62374),
    .lcout(net_58457),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_3 (
    .carryin(net_62370),
    .carryout(net_62376),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62378),
    .in2(net_62379_cascademuxed),
    .in3(net_62380),
    .lcout(net_58458),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_4 (
    .carryin(net_62376),
    .carryout(net_62382),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62384),
    .in2(net_62385_cascademuxed),
    .in3(net_62386),
    .lcout(net_58459),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_5 (
    .carryin(net_62382),
    .carryout(net_62388),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62390),
    .in2(net_62391_cascademuxed),
    .in3(net_62392),
    .lcout(net_58460),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_6 (
    .carryin(net_62388),
    .carryout(net_62394),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62396),
    .in2(net_62397_cascademuxed),
    .in3(net_62398),
    .lcout(net_58461),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_7 (
    .carryin(net_62394),
    .carryout(net_62400),
    .ce(),
    .clk(net_62406),
    .in0(gnd),
    .in1(net_62402),
    .in2(net_62403_cascademuxed),
    .in3(net_62404),
    .lcout(net_58462),
    .ltout(),
    .sr(net_62407)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_17_0 (
    .carryin(net_62444),
    .carryout(net_62481),
    .ce(),
    .clk(net_62529),
    .in0(gnd),
    .in1(net_62483),
    .in2(net_62484_cascademuxed),
    .in3(net_62485),
    .lcout(net_58578),
    .ltout(),
    .sr(net_62530)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_1 (
    .carryin(net_62481),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62491),
    .lcout(net_58579),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62496_cascademuxed),
    .in3(gnd),
    .lcout(net_58580),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_62529),
    .in0(net_62506),
    .in1(net_62507),
    .in2(gnd),
    .in3(net_62509),
    .lcout(net_58582),
    .ltout(),
    .sr(net_62530)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62651),
    .clk(net_62652),
    .in0(net_62629),
    .in1(net_62630),
    .in2(net_62631_cascademuxed),
    .in3(net_62632),
    .lcout(net_58705),
    .ltout(),
    .sr(net_62653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_60683),
    .clk(net_60684),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_60676),
    .lcout(net_56703),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60807),
    .in0(gnd),
    .in1(gnd),
    .in2(net_60774_cascademuxed),
    .in3(gnd),
    .lcout(net_56858),
    .ltout(),
    .sr(net_60808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60807),
    .in0(net_60784),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_56860),
    .ltout(),
    .sr(net_60808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_60886),
    .lcout(net_56979),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(net_60890),
    .in2(gnd),
    .in3(net_60892),
    .lcout(net_56980),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(net_60895),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_56981),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(net_60901),
    .in1(gnd),
    .in2(gnd),
    .in3(net_60904),
    .lcout(net_56982),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(net_60908),
    .in2(net_60909_cascademuxed),
    .in3(gnd),
    .lcout(net_56983),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(net_60914),
    .in2(net_60915_cascademuxed),
    .in3(gnd),
    .lcout(net_56984),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(gnd),
    .in2(net_60921_cascademuxed),
    .in3(net_60922),
    .lcout(net_56985),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_60930),
    .in0(gnd),
    .in1(net_60926),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_56986),
    .ltout(),
    .sr(net_60931)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(net_61006),
    .in1(net_61007),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57102),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(gnd),
    .in1(net_61013),
    .in2(gnd),
    .in3(net_61015),
    .lcout(net_57103),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(net_61018),
    .in1(gnd),
    .in2(net_61020_cascademuxed),
    .in3(gnd),
    .lcout(net_57104),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(gnd),
    .in1(net_61025),
    .in2(gnd),
    .in3(net_61027),
    .lcout(net_57105),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61032_cascademuxed),
    .in3(net_61033),
    .lcout(net_57106),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(net_61036),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61039),
    .lcout(net_57107),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(net_61042),
    .in1(gnd),
    .in2(net_61044_cascademuxed),
    .in3(gnd),
    .lcout(net_57108),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61053),
    .in0(gnd),
    .in1(net_61049),
    .in2(gnd),
    .in3(net_61051),
    .lcout(net_57109),
    .ltout(),
    .sr(net_61054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000011001010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61129),
    .in1(net_61130),
    .in2(net_61131_cascademuxed),
    .in3(net_61132),
    .lcout(net_57225),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61135),
    .in1(net_61136),
    .in2(net_61137_cascademuxed),
    .in3(net_61138),
    .lcout(net_57226),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100101111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61147),
    .in1(net_61148),
    .in2(net_61149_cascademuxed),
    .in3(net_61150),
    .lcout(net_57228),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61153),
    .in1(net_61154),
    .in2(net_61155_cascademuxed),
    .in3(net_61156),
    .lcout(net_57229),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61159),
    .in1(net_61160),
    .in2(net_61161_cascademuxed),
    .in3(net_61162),
    .lcout(net_57230),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61165),
    .in1(net_61166),
    .in2(net_61167_cascademuxed),
    .in3(net_61168),
    .lcout(net_57231),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110010011000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(net_61171),
    .in1(net_61172),
    .in2(net_61173_cascademuxed),
    .in3(net_61174),
    .lcout(net_57232),
    .ltout(),
    .sr(net_61177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61266_cascademuxed),
    .in3(gnd),
    .lcout(net_57350),
    .ltout(),
    .sr(net_61300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61272_cascademuxed),
    .in3(gnd),
    .lcout(net_57351),
    .ltout(),
    .sr(net_61300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61299),
    .in0(net_61276),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57352),
    .ltout(),
    .sr(net_61300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61290_cascademuxed),
    .in3(gnd),
    .lcout(net_57354),
    .ltout(),
    .sr(net_61300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57471),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61422),
    .in0(gnd),
    .in1(net_61382),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57472),
    .ltout(),
    .sr(net_61423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61422),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61390),
    .lcout(net_57473),
    .ltout(),
    .sr(net_61423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61422),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61395_cascademuxed),
    .in3(gnd),
    .lcout(net_57474),
    .ltout(),
    .sr(net_61423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_61422),
    .in0(gnd),
    .in1(net_61400),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57475),
    .ltout(),
    .sr(net_61423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(net_61498),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57594),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61506_cascademuxed),
    .in3(gnd),
    .lcout(net_57595),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61513),
    .lcout(net_57596),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61519),
    .lcout(net_57597),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61524_cascademuxed),
    .in3(gnd),
    .lcout(net_57598),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61536_cascademuxed),
    .in3(gnd),
    .lcout(net_57600),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65454_cascademuxed),
    .in3(net_65455),
    .lcout(net_61547),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65458),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65461),
    .lcout(net_61548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(net_65464),
    .in1(net_65465),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61549),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(net_65470),
    .in1(gnd),
    .in2(net_65472_cascademuxed),
    .in3(gnd),
    .lcout(net_61550),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(gnd),
    .in1(net_65477),
    .in2(net_65478_cascademuxed),
    .in3(gnd),
    .lcout(net_61551),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(net_65482),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65485),
    .lcout(net_61552),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(gnd),
    .in1(net_65489),
    .in2(gnd),
    .in3(net_65491),
    .lcout(net_61553),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65499),
    .in0(net_65494),
    .in1(net_65495),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61554),
    .ltout(),
    .sr(net_65500)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_11_0 (
    .carryin(t853),
    .carryout(net_65574),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65576),
    .in2(net_65577_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_1 (
    .carryin(net_65574),
    .carryout(net_65580),
    .ce(net_65621),
    .clk(net_65622),
    .in0(net_65581),
    .in1(net_65582),
    .in2(net_65583_cascademuxed),
    .in3(net_65584),
    .lcout(net_61671),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_2 (
    .carryin(net_65580),
    .carryout(net_65586),
    .ce(net_65621),
    .clk(net_65622),
    .in0(net_65587),
    .in1(net_65588),
    .in2(net_65589_cascademuxed),
    .in3(net_65590),
    .lcout(net_61672),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_3 (
    .carryin(net_65586),
    .carryout(net_65592),
    .ce(net_65621),
    .clk(net_65622),
    .in0(net_65593),
    .in1(net_65594),
    .in2(net_65595_cascademuxed),
    .in3(net_65596),
    .lcout(net_61673),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_4 (
    .carryin(net_65592),
    .carryout(net_65598),
    .ce(net_65621),
    .clk(net_65622),
    .in0(net_65599),
    .in1(net_65600),
    .in2(net_65601_cascademuxed),
    .in3(net_65602),
    .lcout(net_61674),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_11_5 (
    .carryin(net_65598),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65608),
    .lcout(net_61675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110000001100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65621),
    .clk(net_65622),
    .in0(net_65611),
    .in1(net_65612),
    .in2(net_65613_cascademuxed),
    .in3(gnd),
    .lcout(net_61676),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65621),
    .clk(net_65622),
    .in0(gnd),
    .in1(net_65618),
    .in2(gnd),
    .in3(net_65620),
    .lcout(net_61677),
    .ltout(),
    .sr(net_65623)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65744),
    .clk(net_65745),
    .in0(net_65710),
    .in1(net_65711),
    .in2(net_65712_cascademuxed),
    .in3(net_65713),
    .lcout(net_61795),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65744),
    .clk(net_65745),
    .in0(net_65716),
    .in1(net_65717),
    .in2(net_65718_cascademuxed),
    .in3(net_65719),
    .lcout(net_61796),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010111100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65744),
    .clk(net_65745),
    .in0(net_65734),
    .in1(net_65735),
    .in2(net_65736_cascademuxed),
    .in3(net_65737),
    .lcout(net_61799),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001111100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65744),
    .clk(net_65745),
    .in0(net_65740),
    .in1(net_65741),
    .in2(net_65742_cascademuxed),
    .in3(net_65743),
    .lcout(net_61800),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_0 (
    .carryin(t862),
    .carryout(net_65820),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65822),
    .in2(net_65823_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_1 (
    .carryin(net_65820),
    .carryout(net_65826),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65828),
    .in2(net_65829_cascademuxed),
    .in3(net_65830),
    .lcout(net_61917),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_2 (
    .carryin(net_65826),
    .carryout(net_65832),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65834),
    .in2(net_65835_cascademuxed),
    .in3(net_65836),
    .lcout(net_61918),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_3 (
    .carryin(net_65832),
    .carryout(net_65838),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65840),
    .in2(net_65841_cascademuxed),
    .in3(net_65842),
    .lcout(net_61919),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_4 (
    .carryin(net_65838),
    .carryout(net_65844),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65846),
    .in2(net_65847_cascademuxed),
    .in3(net_65848),
    .lcout(net_61920),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_5 (
    .carryin(net_65844),
    .carryout(net_65850),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65852),
    .in2(net_65853_cascademuxed),
    .in3(net_65854),
    .lcout(net_61921),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_6 (
    .carryin(net_65850),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65860),
    .lcout(net_61922),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65867),
    .clk(net_65868),
    .in0(gnd),
    .in1(net_65864),
    .in2(gnd),
    .in3(net_65866),
    .lcout(net_61923),
    .ltout(),
    .sr(net_65869)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_0 (
    .carryin(t867),
    .carryout(net_65943),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65945),
    .in2(net_65946_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_1 (
    .carryin(net_65943),
    .carryout(net_65949),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65951),
    .in2(net_65952_cascademuxed),
    .in3(net_65953),
    .lcout(net_62040),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_2 (
    .carryin(net_65949),
    .carryout(net_65955),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65957),
    .in2(net_65958_cascademuxed),
    .in3(net_65959),
    .lcout(net_62041),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_3 (
    .carryin(net_65955),
    .carryout(net_65961),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65963),
    .in2(net_65964_cascademuxed),
    .in3(net_65965),
    .lcout(net_62042),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_4 (
    .carryin(net_65961),
    .carryout(net_65967),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65969),
    .in2(net_65970_cascademuxed),
    .in3(net_65971),
    .lcout(net_62043),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_5 (
    .carryin(net_65967),
    .carryout(net_65973),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65975),
    .in2(net_65976_cascademuxed),
    .in3(net_65977),
    .lcout(net_62044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_6 (
    .carryin(net_65973),
    .carryout(net_65979),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65981),
    .in2(net_65982_cascademuxed),
    .in3(net_65983),
    .lcout(net_62045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_7 (
    .carryin(net_65979),
    .carryout(net_65985),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65987),
    .in2(net_65988_cascademuxed),
    .in3(net_65989),
    .lcout(net_62046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001011001101001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66067),
    .in1(gnd),
    .in2(net_66069_cascademuxed),
    .in3(net_66070),
    .lcout(net_62162),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66075_cascademuxed),
    .in3(gnd),
    .lcout(net_62163),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_66080),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62164),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_66114),
    .in0(gnd),
    .in1(net_66086),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62165),
    .ltout(),
    .sr(net_66115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_66114),
    .in0(gnd),
    .in1(net_66092),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62166),
    .ltout(),
    .sr(net_66115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_66114),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_66100),
    .lcout(net_62167),
    .ltout(),
    .sr(net_66115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_66114),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66105_cascademuxed),
    .in3(gnd),
    .lcout(net_62168),
    .ltout(),
    .sr(net_66115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_66112),
    .lcout(net_62169),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110000001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(net_66190),
    .in1(net_66191),
    .in2(net_66192_cascademuxed),
    .in3(net_66193),
    .lcout(net_62285),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(net_66196),
    .in1(net_66197),
    .in2(net_66198_cascademuxed),
    .in3(net_66199),
    .lcout(net_62286),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110000001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(net_66202),
    .in1(net_66203),
    .in2(net_66204_cascademuxed),
    .in3(net_66205),
    .lcout(net_62287),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(gnd),
    .in1(net_66209),
    .in2(net_66210_cascademuxed),
    .in3(gnd),
    .lcout(net_62288),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(gnd),
    .in1(net_66215),
    .in2(net_66216_cascademuxed),
    .in3(gnd),
    .lcout(net_62289),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(gnd),
    .in1(net_66221),
    .in2(gnd),
    .in3(net_66223),
    .lcout(net_62290),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000101010000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(net_66226),
    .in1(net_66227),
    .in2(net_66228_cascademuxed),
    .in3(net_66229),
    .lcout(net_62291),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66234_cascademuxed),
    .in3(net_66235),
    .lcout(net_62292),
    .ltout(),
    .sr(net_66238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(gnd),
    .in1(net_66314),
    .in2(net_66315_cascademuxed),
    .in3(gnd),
    .lcout(net_62408),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66319),
    .in1(gnd),
    .in2(net_66321_cascademuxed),
    .in3(gnd),
    .lcout(net_62409),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66325),
    .in1(net_66326),
    .in2(net_66327_cascademuxed),
    .in3(net_66328),
    .lcout(net_62410),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66331),
    .in1(net_66332),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62411),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(gnd),
    .in1(net_66338),
    .in2(gnd),
    .in3(net_66340),
    .lcout(net_62412),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66343),
    .in1(gnd),
    .in2(net_66345_cascademuxed),
    .in3(gnd),
    .lcout(net_62413),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66349),
    .in1(net_66350),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62414),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(net_66355),
    .in1(net_66356),
    .in2(net_66357_cascademuxed),
    .in3(net_66358),
    .lcout(net_62415),
    .ltout(),
    .sr(net_66361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66482),
    .clk(net_66483),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66438_cascademuxed),
    .in3(gnd),
    .lcout(net_62531),
    .ltout(),
    .sr(net_66484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_64514),
    .clk(net_64515),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64488_cascademuxed),
    .in3(gnd),
    .lcout(net_60530),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111110001111),
    .SEQ_MODE(4'b1000)
  ) lc40_16_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_64637),
    .clk(net_64638),
    .in0(net_64603),
    .in1(net_64604),
    .in2(net_64605_cascademuxed),
    .in3(net_64606),
    .lcout(net_60688),
    .ltout(),
    .sr(net_64639)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111001100),
    .SEQ_MODE(4'b0000)
  ) lc40_16_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64610),
    .in2(gnd),
    .in3(net_64612),
    .lcout(net_60689),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_0 (
    .carryin(t826),
    .carryout(net_64713),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64715),
    .in2(net_64716_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_1 (
    .carryin(net_64713),
    .carryout(net_64719),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64721),
    .in2(net_64722_cascademuxed),
    .in3(net_64723),
    .lcout(net_60810),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_2 (
    .carryin(net_64719),
    .carryout(net_64725),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64727),
    .in2(net_64728_cascademuxed),
    .in3(net_64729),
    .lcout(net_60811),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_3 (
    .carryin(net_64725),
    .carryout(net_64731),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64733),
    .in2(net_64734_cascademuxed),
    .in3(net_64735),
    .lcout(net_60812),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_4 (
    .carryin(net_64731),
    .carryout(net_64737),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64739),
    .in2(net_64740_cascademuxed),
    .in3(net_64741),
    .lcout(net_60813),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_5 (
    .carryin(net_64737),
    .carryout(net_64743),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64745),
    .in2(net_64746_cascademuxed),
    .in3(net_64747),
    .lcout(net_60814),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_6 (
    .carryin(net_64743),
    .carryout(net_64749),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64751),
    .in2(net_64752_cascademuxed),
    .in3(net_64753),
    .lcout(net_60815),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_7 (
    .carryin(net_64749),
    .carryout(net_64755),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64757),
    .in2(net_64758_cascademuxed),
    .in3(net_64759),
    .lcout(net_60816),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_0 (
    .carryin(net_64799),
    .carryout(net_64836),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64838),
    .in2(net_64839_cascademuxed),
    .in3(net_64840),
    .lcout(net_60932),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_1 (
    .carryin(net_64836),
    .carryout(net_64842),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64844),
    .in2(net_64845_cascademuxed),
    .in3(net_64846),
    .lcout(net_60933),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_2 (
    .carryin(net_64842),
    .carryout(net_64848),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64850),
    .in2(net_64851_cascademuxed),
    .in3(net_64852),
    .lcout(net_60934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_3 (
    .carryin(net_64848),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_64858),
    .lcout(net_60935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_64884),
    .in0(net_64861),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_60936),
    .ltout(),
    .sr(net_64885)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64868),
    .in2(gnd),
    .in3(net_64870),
    .lcout(net_60937),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_64884),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_64876),
    .lcout(net_60938),
    .ltout(),
    .sr(net_64885)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_64884),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64881_cascademuxed),
    .in3(gnd),
    .lcout(net_60939),
    .ltout(),
    .sr(net_64885)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_6_0 (
    .carryin(t835),
    .carryout(net_64959),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64961),
    .in2(net_64962_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_1 (
    .carryin(net_64959),
    .carryout(net_64965),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64968_cascademuxed),
    .in3(net_64969),
    .lcout(net_61056),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_2 (
    .carryin(net_64965),
    .carryout(net_64971),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64974_cascademuxed),
    .in3(net_64975),
    .lcout(net_61057),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_3 (
    .carryin(net_64971),
    .carryout(net_64977),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(net_64979),
    .in2(gnd),
    .in3(net_64981),
    .lcout(net_61058),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_4 (
    .carryin(net_64977),
    .carryout(net_64983),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64986_cascademuxed),
    .in3(net_64987),
    .lcout(net_61059),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_5 (
    .carryin(net_64983),
    .carryout(net_64989),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(net_64991),
    .in2(gnd),
    .in3(net_64993),
    .lcout(net_61060),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_6 (
    .carryin(net_64989),
    .carryout(net_64995),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64998_cascademuxed),
    .in3(net_64999),
    .lcout(net_61061),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_6_7 (
    .carryin(net_64995),
    .carryout(net_65001),
    .ce(),
    .clk(net_65007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65004_cascademuxed),
    .in3(net_65005),
    .lcout(net_61062),
    .ltout(),
    .sr(net_65008)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_0 (
    .carryin(net_65045),
    .carryout(net_65082),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65085_cascademuxed),
    .in3(net_65086),
    .lcout(net_61178),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_1 (
    .carryin(net_65082),
    .carryout(net_65088),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(net_65090),
    .in2(gnd),
    .in3(net_65092),
    .lcout(net_61179),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_2 (
    .carryin(net_65088),
    .carryout(net_65094),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(net_65096),
    .in2(gnd),
    .in3(net_65098),
    .lcout(net_61180),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_3 (
    .carryin(net_65094),
    .carryout(net_65100),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65103_cascademuxed),
    .in3(net_65104),
    .lcout(net_61181),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_7_4 (
    .carryin(net_65100),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65110),
    .lcout(net_61182),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65116),
    .lcout(net_61183),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65121_cascademuxed),
    .in3(net_65122),
    .lcout(net_61184),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65130),
    .in0(gnd),
    .in1(net_65126),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61185),
    .ltout(),
    .sr(net_65131)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65253),
    .in0(gnd),
    .in1(net_65207),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61301),
    .ltout(),
    .sr(net_65254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_16_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65253),
    .in0(net_65212),
    .in1(gnd),
    .in2(net_65214_cascademuxed),
    .in3(gnd),
    .lcout(net_61302),
    .ltout(),
    .sr(net_65254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65253),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65232_cascademuxed),
    .in3(gnd),
    .lcout(net_61305),
    .ltout(),
    .sr(net_65254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65337_cascademuxed),
    .in3(gnd),
    .lcout(net_61425),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65344),
    .lcout(net_61426),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65356),
    .lcout(net_61428),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65362),
    .lcout(net_61429),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(net_65366),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61430),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65376),
    .in0(gnd),
    .in1(net_65372),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61431),
    .ltout(),
    .sr(net_65377)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69286),
    .lcout(net_65378),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69292),
    .lcout(net_65379),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(net_69295),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65380),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69303_cascademuxed),
    .in3(gnd),
    .lcout(net_65381),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(net_69308),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65382),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69316),
    .lcout(net_65383),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69330),
    .in0(gnd),
    .in1(net_69326),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65385),
    .ltout(),
    .sr(net_69331)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_0 (
    .carryin(t917),
    .carryout(net_69405),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69407),
    .in2(net_69408_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_1 (
    .carryin(net_69405),
    .carryout(net_69411),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69413),
    .in2(net_69414_cascademuxed),
    .in3(net_69415),
    .lcout(net_65502),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_2 (
    .carryin(net_69411),
    .carryout(net_69417),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69419),
    .in2(net_69420_cascademuxed),
    .in3(net_69421),
    .lcout(net_65503),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_3 (
    .carryin(net_69417),
    .carryout(net_69423),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69425),
    .in2(net_69426_cascademuxed),
    .in3(net_69427),
    .lcout(net_65504),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_4 (
    .carryin(net_69423),
    .carryout(net_69429),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69431),
    .in2(gnd),
    .in3(net_69433),
    .lcout(net_65505),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69436),
    .in1(net_69437),
    .in2(net_69438_cascademuxed),
    .in3(net_69439),
    .lcout(net_65506),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69452),
    .clk(net_69453),
    .in0(net_69442),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69445),
    .lcout(net_65507),
    .ltout(),
    .sr(net_69454)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69452),
    .clk(net_69453),
    .in0(net_69448),
    .in1(net_69449),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65508),
    .ltout(),
    .sr(net_69454)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69532),
    .lcout(net_65624),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(net_69535),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65625),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(net_69541),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65626),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69549_cascademuxed),
    .in3(gnd),
    .lcout(net_65627),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69555_cascademuxed),
    .in3(gnd),
    .lcout(net_65628),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(net_69560),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65629),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69568),
    .lcout(net_65630),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69574),
    .lcout(net_65631),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_0 (
    .carryin(t929),
    .carryout(net_69651),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69653),
    .in2(net_69654_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_1 (
    .carryin(net_69651),
    .carryout(net_69657),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69659),
    .in2(net_69660_cascademuxed),
    .in3(net_69661),
    .lcout(net_65748),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_2 (
    .carryin(net_69657),
    .carryout(net_69663),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69665),
    .in2(net_69666_cascademuxed),
    .in3(net_69667),
    .lcout(net_65749),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_3 (
    .carryin(net_69663),
    .carryout(net_69669),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69671),
    .in2(net_69672_cascademuxed),
    .in3(net_69673),
    .lcout(net_65750),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_4 (
    .carryin(net_69669),
    .carryout(net_69675),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69677),
    .in2(net_69678_cascademuxed),
    .in3(net_69679),
    .lcout(net_65751),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_5 (
    .carryin(net_69675),
    .carryout(net_69681),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69683),
    .in2(net_69684_cascademuxed),
    .in3(net_69685),
    .lcout(net_65752),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_6 (
    .carryin(net_69681),
    .carryout(t1004),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69689),
    .in2(net_69690_cascademuxed),
    .in3(net_69691),
    .lcout(net_65753),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_13_7 (
    .carryin(t1004),
    .carryout(net_69693),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_69695),
    .in2(net_69696_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69775),
    .in1(gnd),
    .in2(net_69777_cascademuxed),
    .in3(net_69778),
    .lcout(net_65870),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69821),
    .clk(net_69822),
    .in0(net_69781),
    .in1(net_69782),
    .in2(net_69783_cascademuxed),
    .in3(net_69784),
    .lcout(net_65871),
    .ltout(),
    .sr(net_69823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100100000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69821),
    .clk(net_69822),
    .in0(net_69787),
    .in1(net_69788),
    .in2(net_69789_cascademuxed),
    .in3(net_69790),
    .lcout(net_65872),
    .ltout(),
    .sr(net_69823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110000001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69821),
    .clk(net_69822),
    .in0(net_69793),
    .in1(net_69794),
    .in2(net_69795_cascademuxed),
    .in3(net_69796),
    .lcout(net_65873),
    .ltout(),
    .sr(net_69823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69799),
    .in1(net_69800),
    .in2(net_69801_cascademuxed),
    .in3(gnd),
    .lcout(net_65874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_17_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69808),
    .lcout(net_65875),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100100001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69821),
    .clk(net_69822),
    .in0(net_69811),
    .in1(net_69812),
    .in2(net_69813_cascademuxed),
    .in3(net_69814),
    .lcout(net_65876),
    .ltout(),
    .sr(net_69823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69821),
    .clk(net_69822),
    .in0(net_69817),
    .in1(net_69818),
    .in2(net_69819_cascademuxed),
    .in3(net_69820),
    .lcout(net_65877),
    .ltout(),
    .sr(net_69823)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_17_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69900_cascademuxed),
    .in3(gnd),
    .lcout(net_65993),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(gnd),
    .in1(net_69905),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65994),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(gnd),
    .in1(net_69911),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65995),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_17_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69918_cascademuxed),
    .in3(gnd),
    .lcout(net_65996),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69925),
    .lcout(net_65997),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(gnd),
    .in1(gnd),
    .in2(net_69930_cascademuxed),
    .in3(gnd),
    .lcout(net_65998),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(net_69934),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65999),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69945),
    .in0(net_69940),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66000),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_0 (
    .carryin(t948),
    .carryout(net_70020),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70022),
    .in2(net_70023_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_1 (
    .carryin(net_70020),
    .carryout(net_70026),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70028),
    .in2(gnd),
    .in3(net_70030),
    .lcout(net_66117),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_2 (
    .carryin(net_70026),
    .carryout(net_70032),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70035_cascademuxed),
    .in3(net_70036),
    .lcout(net_66118),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_3 (
    .carryin(net_70032),
    .carryout(net_70038),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70041_cascademuxed),
    .in3(net_70042),
    .lcout(net_66119),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_4 (
    .carryin(net_70038),
    .carryout(net_70044),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70046),
    .in2(gnd),
    .in3(net_70048),
    .lcout(net_66120),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_5 (
    .carryin(net_70044),
    .carryout(net_70050),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70052),
    .in2(gnd),
    .in3(net_70054),
    .lcout(net_66121),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_6 (
    .carryin(net_70050),
    .carryout(t957),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70058),
    .in2(gnd),
    .in3(net_70060),
    .lcout(net_66122),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_7 (
    .carryin(t957),
    .carryout(net_70062),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70064),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_0 (
    .carryin(net_70106),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70147),
    .lcout(net_66239),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010100000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(net_70150),
    .in1(net_70151),
    .in2(net_70152_cascademuxed),
    .in3(net_70153),
    .lcout(net_66240),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70163),
    .in2(gnd),
    .in3(net_70165),
    .lcout(net_66242),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(net_70168),
    .in1(net_70169),
    .in2(net_70170_cascademuxed),
    .in3(net_70171),
    .lcout(net_66243),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70174),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70177),
    .lcout(net_66244),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000110010000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(net_70180),
    .in1(net_70181),
    .in2(net_70182_cascademuxed),
    .in3(net_70183),
    .lcout(net_66245),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(net_70186),
    .in1(net_70187),
    .in2(net_70188_cascademuxed),
    .in3(net_70189),
    .lcout(net_66246),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(net_70303),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66368),
    .ltout(),
    .sr(net_70315)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68345),
    .clk(net_68346),
    .in0(net_68299),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64358),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68345),
    .clk(net_68346),
    .in0(net_68341),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64365),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68424_cascademuxed),
    .in3(gnd),
    .lcout(net_64517),
    .ltout(),
    .sr(net_68470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68430_cascademuxed),
    .in3(gnd),
    .lcout(net_64518),
    .ltout(),
    .sr(net_68470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68436_cascademuxed),
    .in3(gnd),
    .lcout(net_64519),
    .ltout(),
    .sr(net_68470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68469),
    .in0(net_68440),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64520),
    .ltout(),
    .sr(net_68470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68469),
    .in0(net_68446),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64521),
    .ltout(),
    .sr(net_68470)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(net_68546),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64640),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68553_cascademuxed),
    .in3(gnd),
    .lcout(net_64641),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_68560),
    .lcout(net_64642),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_68566),
    .lcout(net_64643),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_68572),
    .lcout(net_64644),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_68578),
    .lcout(net_64645),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68583_cascademuxed),
    .in3(gnd),
    .lcout(net_64646),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68592),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68589_cascademuxed),
    .in3(gnd),
    .lcout(net_64647),
    .ltout(),
    .sr(net_68593)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68670_cascademuxed),
    .in3(gnd),
    .lcout(net_64763),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(net_68674),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64764),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68682_cascademuxed),
    .in3(gnd),
    .lcout(net_64765),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(gnd),
    .in1(net_68687),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64766),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(net_68698),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64768),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68706_cascademuxed),
    .in3(gnd),
    .lcout(net_64769),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68712_cascademuxed),
    .in3(gnd),
    .lcout(net_64770),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68838),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68805_cascademuxed),
    .in3(gnd),
    .lcout(net_64888),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68838),
    .in0(net_68815),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64890),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68838),
    .in0(gnd),
    .in1(net_68822),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64891),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68838),
    .in0(net_68827),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64892),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_68838),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68835_cascademuxed),
    .in3(gnd),
    .lcout(net_64893),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b1000)
  ) lc40_17_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68960),
    .clk(net_68961),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68958_cascademuxed),
    .in3(gnd),
    .lcout(net_65016),
    .ltout(),
    .sr(net_68962)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011011000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69083),
    .clk(net_69084),
    .in0(net_69043),
    .in1(net_69044),
    .in2(net_69045_cascademuxed),
    .in3(net_69046),
    .lcout(net_65133),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69083),
    .clk(net_69084),
    .in0(net_69049),
    .in1(net_69050),
    .in2(net_69051_cascademuxed),
    .in3(net_69052),
    .lcout(net_65134),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69083),
    .clk(net_69084),
    .in0(net_69073),
    .in1(net_69074),
    .in2(net_69075_cascademuxed),
    .in3(net_69076),
    .lcout(net_65138),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69207),
    .in0(gnd),
    .in1(net_69185),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65259),
    .ltout(),
    .sr(net_69208)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69207),
    .in0(gnd),
    .in1(net_69203),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65262),
    .ltout(),
    .sr(net_69208)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_10_0 (
    .carryin(t987),
    .carryout(net_73113),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73115),
    .in2(net_73116_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_1 (
    .carryin(net_73113),
    .carryout(net_73119),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73121),
    .in2(net_73122_cascademuxed),
    .in3(net_73123),
    .lcout(net_69210),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_2 (
    .carryin(net_73119),
    .carryout(net_73125),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73127),
    .in2(net_73128_cascademuxed),
    .in3(net_73129),
    .lcout(net_69211),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_3 (
    .carryin(net_73125),
    .carryout(net_73131),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73133),
    .in2(net_73134_cascademuxed),
    .in3(net_73135),
    .lcout(net_69212),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_4 (
    .carryin(net_73131),
    .carryout(net_73137),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73139),
    .in2(net_73140_cascademuxed),
    .in3(net_73141),
    .lcout(net_69213),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_5 (
    .carryin(net_73137),
    .carryout(net_73143),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73145),
    .in2(net_73146_cascademuxed),
    .in3(net_73147),
    .lcout(net_69214),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_10_6 (
    .carryin(net_73143),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73153),
    .lcout(net_69215),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73161),
    .in0(gnd),
    .in1(net_73157),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69216),
    .ltout(),
    .sr(net_73162)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73240),
    .lcout(net_69332),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(net_73243),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69333),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(gnd),
    .in1(net_73250),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69334),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73258),
    .lcout(net_69335),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73264),
    .lcout(net_69336),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(net_73267),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69337),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73275_cascademuxed),
    .in3(gnd),
    .lcout(net_69338),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73284),
    .in0(net_73279),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69339),
    .ltout(),
    .sr(net_73285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(net_73360),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69455),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(net_73367),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69456),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73375),
    .lcout(net_69457),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73381),
    .lcout(net_69458),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73386_cascademuxed),
    .in3(gnd),
    .lcout(net_69459),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73399),
    .lcout(net_69461),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73404_cascademuxed),
    .in3(gnd),
    .lcout(net_69462),
    .ltout(),
    .sr(net_73408)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73486),
    .lcout(net_69578),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73492),
    .lcout(net_69579),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73497_cascademuxed),
    .in3(gnd),
    .lcout(net_69580),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(net_73507),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69582),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(net_73513),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69583),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73521_cascademuxed),
    .in3(gnd),
    .lcout(net_69584),
    .ltout(),
    .sr(net_73531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73608_cascademuxed),
    .in3(gnd),
    .lcout(net_69701),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(net_73612),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69702),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(net_73618),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69703),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73626_cascademuxed),
    .in3(gnd),
    .lcout(net_69704),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(net_73631),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69705),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(net_73637),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69706),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(net_73643),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69707),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73653),
    .in0(gnd),
    .in1(net_73649),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69708),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_0 (
    .carryin(t1013),
    .carryout(net_73728),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73730),
    .in2(net_73731_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_1 (
    .carryin(net_73728),
    .carryout(net_73734),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73736),
    .in2(net_73737_cascademuxed),
    .in3(net_73738),
    .lcout(net_69825),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_2 (
    .carryin(net_73734),
    .carryout(net_73740),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73742),
    .in2(net_73743_cascademuxed),
    .in3(net_73744),
    .lcout(net_69826),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_3 (
    .carryin(net_73740),
    .carryout(net_73746),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73748),
    .in2(net_73749_cascademuxed),
    .in3(net_73750),
    .lcout(net_69827),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_4 (
    .carryin(net_73746),
    .carryout(net_73752),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73754),
    .in2(net_73755_cascademuxed),
    .in3(net_73756),
    .lcout(net_69828),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_5 (
    .carryin(net_73752),
    .carryout(net_73758),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73760),
    .in2(net_73761_cascademuxed),
    .in3(net_73762),
    .lcout(net_69829),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_6 (
    .carryin(net_73758),
    .carryout(net_73764),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73766),
    .in2(net_73767_cascademuxed),
    .in3(net_73768),
    .lcout(net_69830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_15_7 (
    .carryin(net_73764),
    .carryout(net_73770),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73772),
    .in2(net_73773_cascademuxed),
    .in3(net_73774),
    .lcout(net_69831),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73852),
    .in1(net_73853),
    .in2(net_73854_cascademuxed),
    .in3(net_73855),
    .lcout(net_69947),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73899),
    .in0(gnd),
    .in1(net_73859),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69948),
    .ltout(),
    .sr(net_73900)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73899),
    .in0(net_73864),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69949),
    .ltout(),
    .sr(net_73900)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73876),
    .in1(gnd),
    .in2(net_73878_cascademuxed),
    .in3(gnd),
    .lcout(net_69951),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73899),
    .in0(gnd),
    .in1(net_73883),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69952),
    .ltout(),
    .sr(net_73900)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73899),
    .in0(gnd),
    .in1(net_73895),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69954),
    .ltout(),
    .sr(net_73900)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(net_73999),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70074),
    .ltout(),
    .sr(net_74023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72177),
    .in0(net_72154),
    .in1(net_72155),
    .in2(gnd),
    .in3(net_72157),
    .lcout(net_68193),
    .ltout(),
    .sr(net_72178)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(net_72253),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68348),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72261_cascademuxed),
    .in3(gnd),
    .lcout(net_68349),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72267_cascademuxed),
    .in3(gnd),
    .lcout(net_68350),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(net_72272),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68351),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72279_cascademuxed),
    .in3(gnd),
    .lcout(net_68352),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72285_cascademuxed),
    .in3(gnd),
    .lcout(net_68353),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(net_72289),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68354),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72300),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72298),
    .lcout(net_68355),
    .ltout(),
    .sr(net_72301)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_0 (
    .carryin(t968),
    .carryout(net_72375),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72377),
    .in2(net_72378_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_1 (
    .carryin(net_72375),
    .carryout(net_72381),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72383),
    .in2(net_72384_cascademuxed),
    .in3(net_72385),
    .lcout(net_68472),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_2 (
    .carryin(net_72381),
    .carryout(net_72387),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72389),
    .in2(net_72390_cascademuxed),
    .in3(net_72391),
    .lcout(net_68473),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_3 (
    .carryin(net_72387),
    .carryout(net_72393),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72395),
    .in2(net_72396_cascademuxed),
    .in3(net_72397),
    .lcout(net_68474),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_4 (
    .carryin(net_72393),
    .carryout(net_72399),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72401),
    .in2(net_72402_cascademuxed),
    .in3(net_72403),
    .lcout(net_68475),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_5 (
    .carryin(net_72399),
    .carryout(net_72405),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72407),
    .in2(net_72408_cascademuxed),
    .in3(net_72409),
    .lcout(net_68476),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_6 (
    .carryin(net_72405),
    .carryout(net_72411),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72413),
    .in2(net_72414_cascademuxed),
    .in3(net_72415),
    .lcout(net_68477),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_4_7 (
    .carryin(net_72411),
    .carryout(net_72417),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72419),
    .in2(net_72420_cascademuxed),
    .in3(net_72421),
    .lcout(net_68478),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_5_0 (
    .carryin(net_72461),
    .carryout(net_72498),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72500),
    .in2(net_72501_cascademuxed),
    .in3(net_72502),
    .lcout(net_68594),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72505),
    .in1(net_72506),
    .in2(gnd),
    .in3(net_72508),
    .lcout(net_68595),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(net_72511),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68596),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72520),
    .lcout(net_68597),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(gnd),
    .in1(net_72524),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68598),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72532),
    .lcout(net_68599),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72537_cascademuxed),
    .in3(gnd),
    .lcout(net_68600),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72546),
    .in0(gnd),
    .in1(net_72542),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68601),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72624_cascademuxed),
    .in3(gnd),
    .lcout(net_68717),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72630_cascademuxed),
    .in3(gnd),
    .lcout(net_68718),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(gnd),
    .in1(gnd),
    .in2(net_72642_cascademuxed),
    .in3(gnd),
    .lcout(net_68720),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(gnd),
    .in1(net_72647),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68721),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(net_72652),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68722),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72669),
    .in0(net_72658),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68723),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72664),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72667),
    .lcout(net_68724),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_7_0 (
    .carryin(t980),
    .carryout(net_72744),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72746),
    .in2(net_72747_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_1 (
    .carryin(net_72744),
    .carryout(net_72750),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72752),
    .in2(net_72753_cascademuxed),
    .in3(net_72754),
    .lcout(net_68841),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_2 (
    .carryin(net_72750),
    .carryout(net_72756),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72758),
    .in2(net_72759_cascademuxed),
    .in3(net_72760),
    .lcout(net_68842),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_3 (
    .carryin(net_72756),
    .carryout(net_72762),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72764),
    .in2(net_72765_cascademuxed),
    .in3(net_72766),
    .lcout(net_68843),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_4 (
    .carryin(net_72762),
    .carryout(net_72768),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72770),
    .in2(net_72771_cascademuxed),
    .in3(net_72772),
    .lcout(net_68844),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_5 (
    .carryin(net_72768),
    .carryout(net_72774),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72776),
    .in2(net_72777_cascademuxed),
    .in3(net_72778),
    .lcout(net_68845),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_6 (
    .carryin(net_72774),
    .carryout(net_72780),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72782),
    .in2(net_72783_cascademuxed),
    .in3(net_72784),
    .lcout(net_68846),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_7_7 (
    .carryin(net_72780),
    .carryout(net_72786),
    .ce(),
    .clk(net_72792),
    .in0(gnd),
    .in1(net_72788),
    .in2(net_72789_cascademuxed),
    .in3(net_72790),
    .lcout(net_68847),
    .ltout(),
    .sr(net_72793)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_8_0 (
    .carryin(net_72830),
    .carryout(net_72867),
    .ce(),
    .clk(net_72915),
    .in0(gnd),
    .in1(net_72869),
    .in2(net_72870_cascademuxed),
    .in3(net_72871),
    .lcout(net_68963),
    .ltout(),
    .sr(net_72916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72915),
    .in0(net_72874),
    .in1(net_72875),
    .in2(gnd),
    .in3(net_72877),
    .lcout(net_68964),
    .ltout(),
    .sr(net_72916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72915),
    .in0(gnd),
    .in1(net_72893),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68967),
    .ltout(),
    .sr(net_72916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72915),
    .in0(net_72898),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_68968),
    .ltout(),
    .sr(net_72916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_72915),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72913),
    .lcout(net_68970),
    .ltout(),
    .sr(net_72916)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73038),
    .in0(net_72991),
    .in1(gnd),
    .in2(net_72993_cascademuxed),
    .in3(gnd),
    .lcout(net_69086),
    .ltout(),
    .sr(net_73039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73038),
    .in0(net_72997),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69087),
    .ltout(),
    .sr(net_73039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73038),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73012),
    .lcout(net_69089),
    .ltout(),
    .sr(net_73039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73038),
    .in0(gnd),
    .in1(net_73022),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69091),
    .ltout(),
    .sr(net_73039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73038),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73029_cascademuxed),
    .in3(gnd),
    .lcout(net_69092),
    .ltout(),
    .sr(net_73039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8114),
    .lcout(net_1965),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8120),
    .lcout(net_1966),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(net_8124),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1967),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8131_cascademuxed),
    .in3(gnd),
    .lcout(net_1968),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(net_8136),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1969),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8143_cascademuxed),
    .in3(gnd),
    .lcout(net_1970),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8149_cascademuxed),
    .in3(gnd),
    .lcout(net_1971),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8158),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8155_cascademuxed),
    .in3(gnd),
    .lcout(net_1972),
    .ltout(),
    .sr(net_8159)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8261),
    .lcout(net_2190),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8266_cascademuxed),
    .in3(gnd),
    .lcout(net_2191),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(net_8271),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2192),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(net_8276),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2193),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(net_8283),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2194),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8291),
    .lcout(net_2195),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(net_8294),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2196),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8305),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8303),
    .lcout(net_2197),
    .ltout(),
    .sr(net_8306)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(net_8406),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2396),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(net_8418),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2398),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(net_8424),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2399),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(net_8430),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2400),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8438),
    .lcout(net_2401),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8444),
    .lcout(net_2402),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8452),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8450),
    .lcout(net_2403),
    .ltout(),
    .sr(net_8453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(gnd),
    .in1(net_8553),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2604),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8560_cascademuxed),
    .in3(gnd),
    .lcout(net_2605),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(net_8564),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2606),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8573),
    .lcout(net_2607),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(net_8576),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2608),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(net_8582),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2609),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8591),
    .lcout(net_2610),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8599),
    .in0(net_8594),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2611),
    .ltout(),
    .sr(net_8600)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(net_8700),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2813),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8707_cascademuxed),
    .in3(gnd),
    .lcout(net_2814),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8714),
    .lcout(net_2815),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8719_cascademuxed),
    .in3(gnd),
    .lcout(net_2816),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8726),
    .lcout(net_2817),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(net_8730),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2818),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(net_8735),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_2819),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8746),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8743_cascademuxed),
    .in3(gnd),
    .lcout(net_2820),
    .ltout(),
    .sr(net_8747)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(net_8846),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3025),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8854_cascademuxed),
    .in3(gnd),
    .lcout(net_3026),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8861),
    .lcout(net_3027),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(gnd),
    .in1(gnd),
    .in2(net_8866_cascademuxed),
    .in3(gnd),
    .lcout(net_3028),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(net_8870),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3029),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8879),
    .lcout(net_3030),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(net_8882),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3031),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8893),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8891),
    .lcout(net_3032),
    .ltout(),
    .sr(net_8894)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_8996),
    .lcout(net_3250),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9001_cascademuxed),
    .in3(gnd),
    .lcout(net_3251),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_9008),
    .lcout(net_3252),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_9014),
    .lcout(net_3253),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(net_9018),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3254),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(net_9024),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3255),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9040),
    .in0(gnd),
    .in1(net_9030),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3256),
    .ltout(),
    .sr(net_9041)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9187),
    .in0(net_9146),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3457),
    .ltout(),
    .sr(net_9188)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9187),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9154_cascademuxed),
    .in3(gnd),
    .lcout(net_3458),
    .ltout(),
    .sr(net_9188)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9187),
    .in0(gnd),
    .in1(net_9159),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3459),
    .ltout(),
    .sr(net_9188)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9187),
    .in0(net_9182),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3463),
    .ltout(),
    .sr(net_9188)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9334),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9289_cascademuxed),
    .in3(gnd),
    .lcout(net_3664),
    .ltout(),
    .sr(net_9335)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9334),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9295_cascademuxed),
    .in3(gnd),
    .lcout(net_3665),
    .ltout(),
    .sr(net_9335)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9334),
    .in0(net_9311),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3668),
    .ltout(),
    .sr(net_9335)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9334),
    .in0(net_9323),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3670),
    .ltout(),
    .sr(net_9335)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9481),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9436_cascademuxed),
    .in3(gnd),
    .lcout(net_3873),
    .ltout(),
    .sr(net_9482)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9481),
    .in0(gnd),
    .in1(net_9465),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3878),
    .ltout(),
    .sr(net_9482)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9481),
    .in0(net_9476),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_3880),
    .ltout(),
    .sr(net_9482)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_1_1_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_6760),
    .in1(net_6761),
    .in2(gnd),
    .in3(net_6763),
    .lcout(net_103),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110110001000),
    .SEQ_MODE(4'b0000)
  ) lc40_1_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_6778),
    .in1(net_6779),
    .in2(gnd),
    .in3(net_6781),
    .lcout(net_106),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_6795),
    .in0(net_6784),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_107),
    .ltout(),
    .sr(net_6796)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_6795),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6792_cascademuxed),
    .in3(gnd),
    .lcout(net_108),
    .ltout(),
    .sr(net_6796)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9628),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_9590),
    .lcout(net_4086),
    .ltout(),
    .sr(net_9629)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9628),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_9596),
    .lcout(net_4087),
    .ltout(),
    .sr(net_9629)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_20_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9628),
    .in0(net_9617),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_4091),
    .ltout(),
    .sr(net_9629)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9628),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9625_cascademuxed),
    .in3(gnd),
    .lcout(net_4092),
    .ltout(),
    .sr(net_9629)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_21_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9775),
    .in0(gnd),
    .in1(net_9729),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_4312),
    .ltout(),
    .sr(net_9776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_21_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9775),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9748_cascademuxed),
    .in3(gnd),
    .lcout(net_4315),
    .ltout(),
    .sr(net_9776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_22_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9922),
    .in0(gnd),
    .in1(net_9882),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_4540),
    .ltout(),
    .sr(net_9923)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_22_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9922),
    .in0(net_9905),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_4544),
    .ltout(),
    .sr(net_9923)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_22_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_9922),
    .in0(gnd),
    .in1(gnd),
    .in2(net_9913_cascademuxed),
    .in3(gnd),
    .lcout(net_4545),
    .ltout(),
    .sr(net_9923)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_23_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_10069),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_10037),
    .lcout(net_4768),
    .ltout(),
    .sr(net_10070)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_1_2_0 (
    .carryin(t0),
    .carryout(t2),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6937_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_1 (
    .carryin(t2),
    .carryout(net_6940),
    .ce(),
    .clk(net_6982),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6943_cascademuxed),
    .in3(net_6944),
    .lcout(net_117),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_2 (
    .carryin(net_6940),
    .carryout(net_6946),
    .ce(),
    .clk(net_6982),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6949_cascademuxed),
    .in3(net_6950),
    .lcout(net_118),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_3 (
    .carryin(net_6946),
    .carryout(net_6952),
    .ce(),
    .clk(net_6982),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6955_cascademuxed),
    .in3(net_6956),
    .lcout(net_119),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_4 (
    .carryin(net_6952),
    .carryout(net_6958),
    .ce(),
    .clk(net_6982),
    .in0(gnd),
    .in1(net_6960),
    .in2(gnd),
    .in3(net_6962),
    .lcout(net_120),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_5 (
    .carryin(net_6958),
    .carryout(net_6964),
    .ce(),
    .clk(net_6982),
    .in0(gnd),
    .in1(gnd),
    .in2(net_6967_cascademuxed),
    .in3(net_6968),
    .lcout(net_121),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_6982),
    .in0(net_6971),
    .in1(gnd),
    .in2(gnd),
    .in3(net_6974),
    .lcout(net_122),
    .ltout(),
    .sr(net_6983)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001000000001001),
    .SEQ_MODE(4'b0000)
  ) lc40_1_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_6977),
    .in1(net_6978),
    .in2(net_6979_cascademuxed),
    .in3(net_6980),
    .lcout(net_123),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_1_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_7082),
    .in1(gnd),
    .in2(net_7084_cascademuxed),
    .in3(net_7085),
    .lcout(net_451),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011100010),
    .SEQ_MODE(4'b0000)
  ) lc40_1_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_7088),
    .in1(net_7089),
    .in2(net_7090_cascademuxed),
    .in3(gnd),
    .lcout(net_452),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7096_cascademuxed),
    .in3(gnd),
    .lcout(net_453),
    .ltout(),
    .sr(net_7130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7129),
    .in0(net_7100),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_454),
    .ltout(),
    .sr(net_7130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7108_cascademuxed),
    .in3(gnd),
    .lcout(net_455),
    .ltout(),
    .sr(net_7130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7114_cascademuxed),
    .in3(gnd),
    .lcout(net_456),
    .ltout(),
    .sr(net_7130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000100001),
    .SEQ_MODE(4'b0000)
  ) lc40_1_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_7118),
    .in1(net_7119),
    .in2(net_7120_cascademuxed),
    .in3(net_7121),
    .lcout(net_457),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101000001010),
    .SEQ_MODE(4'b0000)
  ) lc40_1_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_7124),
    .in1(gnd),
    .in2(net_7126_cascademuxed),
    .in3(net_7127),
    .lcout(net_458),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_1_4_0 (
    .carryin(t3),
    .carryout(t5),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7231_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_1 (
    .carryin(t5),
    .carryout(net_7234),
    .ce(),
    .clk(net_7276),
    .in0(gnd),
    .in1(net_7236),
    .in2(gnd),
    .in3(net_7238),
    .lcout(net_679),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_2 (
    .carryin(net_7234),
    .carryout(net_7240),
    .ce(),
    .clk(net_7276),
    .in0(gnd),
    .in1(net_7242),
    .in2(gnd),
    .in3(net_7244),
    .lcout(net_680),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_3 (
    .carryin(net_7240),
    .carryout(net_7246),
    .ce(),
    .clk(net_7276),
    .in0(gnd),
    .in1(net_7248),
    .in2(gnd),
    .in3(net_7250),
    .lcout(net_681),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_4 (
    .carryin(net_7246),
    .carryout(net_7252),
    .ce(),
    .clk(net_7276),
    .in0(gnd),
    .in1(net_7254),
    .in2(gnd),
    .in3(net_7256),
    .lcout(net_682),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_5 (
    .carryin(net_7252),
    .carryout(net_7258),
    .ce(),
    .clk(net_7276),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7261_cascademuxed),
    .in3(net_7262),
    .lcout(net_683),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_1_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7276),
    .in0(net_7265),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7268),
    .lcout(net_684),
    .ltout(),
    .sr(net_7277)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000001001000001),
    .SEQ_MODE(4'b0000)
  ) lc40_1_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_7271),
    .in1(net_7272),
    .in2(net_7273_cascademuxed),
    .in3(net_7274),
    .lcout(net_685),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(net_7377),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_905),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7384_cascademuxed),
    .in3(gnd),
    .lcout(net_906),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7390_cascademuxed),
    .in3(gnd),
    .lcout(net_907),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(net_7395),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_908),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7402_cascademuxed),
    .in3(gnd),
    .lcout(net_909),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_1_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_7407),
    .in2(net_7408_cascademuxed),
    .in3(net_7409),
    .lcout(net_910),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7415),
    .lcout(net_911),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7423),
    .in0(net_7418),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_912),
    .ltout(),
    .sr(net_7424)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7570),
    .in0(net_7529),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1131),
    .ltout(),
    .sr(net_7571)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7570),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7543_cascademuxed),
    .in3(gnd),
    .lcout(net_1133),
    .ltout(),
    .sr(net_7571)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7570),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7549_cascademuxed),
    .in3(gnd),
    .lcout(net_1134),
    .ltout(),
    .sr(net_7571)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7570),
    .in0(gnd),
    .in1(net_7554),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1135),
    .ltout(),
    .sr(net_7571)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7570),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7561_cascademuxed),
    .in3(gnd),
    .lcout(net_1136),
    .ltout(),
    .sr(net_7571)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_7716),
    .clk(net_7717),
    .in0(net_7676),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1337),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(net_7817),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1544),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(net_7823),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1545),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7832),
    .lcout(net_1546),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(net_7835),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1547),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(gnd),
    .in1(net_7842),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1548),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7850),
    .lcout(net_1549),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(net_7853),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1550),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_7864),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7861_cascademuxed),
    .in3(gnd),
    .lcout(net_1551),
    .ltout(),
    .sr(net_7865)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(gnd),
    .in1(gnd),
    .in2(net_7966_cascademuxed),
    .in3(gnd),
    .lcout(net_1753),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7973),
    .lcout(net_1754),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(gnd),
    .in1(net_7977),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1755),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(net_7982),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1756),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(net_7988),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1757),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_7997),
    .lcout(net_1758),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(net_8000),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1759),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_1_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_8011),
    .in0(gnd),
    .in1(net_8007),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_1760),
    .ltout(),
    .sr(net_8012)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80191),
    .clk(net_80192),
    .in0(gnd),
    .in1(net_80146),
    .in2(gnd),
    .in3(net_80148),
    .lcout(net_76651),
    .ltout(),
    .sr(net_80193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80191),
    .clk(net_80192),
    .in0(net_80151),
    .in1(net_80152),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76652),
    .ltout(),
    .sr(net_80193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80191),
    .clk(net_80192),
    .in0(net_80169),
    .in1(net_80170),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76655),
    .ltout(),
    .sr(net_80193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80191),
    .clk(net_80192),
    .in0(net_80175),
    .in1(gnd),
    .in2(net_80177_cascademuxed),
    .in3(gnd),
    .lcout(net_76656),
    .ltout(),
    .sr(net_80193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80315),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_80307),
    .lcout(net_76759),
    .ltout(),
    .sr(net_80316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80315),
    .in0(gnd),
    .in1(net_80311),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76760),
    .ltout(),
    .sr(net_80316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(net_80403),
    .in1(gnd),
    .in2(net_80405_cascademuxed),
    .in3(gnd),
    .lcout(net_76857),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80683),
    .clk(net_80684),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_80658),
    .lcout(net_77062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000101),
    .SEQ_MODE(4'b1000)
  ) lc40_20_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79207),
    .clk(net_79208),
    .in0(net_79173),
    .in1(gnd),
    .in2(net_79175_cascademuxed),
    .in3(gnd),
    .lcout(net_75801),
    .ltout(),
    .sr(net_79209)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011001100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79207),
    .clk(net_79208),
    .in0(gnd),
    .in1(net_79204),
    .in2(gnd),
    .in3(net_79206),
    .lcout(net_75806),
    .ltout(),
    .sr(net_79209)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_79287),
    .lcout(net_75937),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_79293),
    .lcout(net_75938),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(net_79302),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_75940),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(net_79314),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_75942),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(net_79320),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_75943),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79331),
    .in0(net_79326),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_75944),
    .ltout(),
    .sr(net_79332)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79453),
    .clk(net_79454),
    .in0(gnd),
    .in1(net_79414),
    .in2(net_79415_cascademuxed),
    .in3(gnd),
    .lcout(net_76040),
    .ltout(),
    .sr(net_79455)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(net_79530),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76141),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(gnd),
    .in2(net_79538_cascademuxed),
    .in3(gnd),
    .lcout(net_76142),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(net_79543),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76143),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_79551),
    .lcout(net_76144),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(net_79554),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76145),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_79563),
    .lcout(net_76146),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_79569),
    .lcout(net_76147),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79577),
    .in0(gnd),
    .in1(net_79573),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76148),
    .ltout(),
    .sr(net_79578)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79699),
    .clk(net_79700),
    .in0(net_79653),
    .in1(net_79654),
    .in2(net_79655_cascademuxed),
    .in3(net_79656),
    .lcout(net_76243),
    .ltout(),
    .sr(net_79701)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79699),
    .clk(net_79700),
    .in0(net_79677),
    .in1(net_79678),
    .in2(net_79679_cascademuxed),
    .in3(net_79680),
    .lcout(net_76247),
    .ltout(),
    .sr(net_79701)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111010100100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79699),
    .clk(net_79700),
    .in0(net_79683),
    .in1(net_79684),
    .in2(net_79685_cascademuxed),
    .in3(net_79686),
    .lcout(net_76248),
    .ltout(),
    .sr(net_79701)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79822),
    .clk(net_79823),
    .in0(net_79806),
    .in1(net_79807),
    .in2(net_79808_cascademuxed),
    .in3(net_79809),
    .lcout(net_76350),
    .ltout(),
    .sr(net_79824)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_79946),
    .in0(gnd),
    .in1(gnd),
    .in2(net_79937_cascademuxed),
    .in3(gnd),
    .lcout(net_76453),
    .ltout(),
    .sr(net_79947)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80069),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_80043),
    .lcout(net_76552),
    .ltout(),
    .sr(net_80070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80069),
    .in0(gnd),
    .in1(gnd),
    .in2(net_80048_cascademuxed),
    .in3(gnd),
    .lcout(net_76553),
    .ltout(),
    .sr(net_80070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80069),
    .in0(gnd),
    .in1(net_80053),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76554),
    .ltout(),
    .sr(net_80070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80069),
    .in0(gnd),
    .in1(gnd),
    .in2(net_80066_cascademuxed),
    .in3(gnd),
    .lcout(net_76556),
    .ltout(),
    .sr(net_80070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84023),
    .in0(net_83976),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80071),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84023),
    .in0(gnd),
    .in1(net_83983),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80072),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84023),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83990_cascademuxed),
    .in3(gnd),
    .lcout(net_80073),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84023),
    .in0(gnd),
    .in1(net_83995),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80074),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84023),
    .in0(gnd),
    .in1(net_84001),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80075),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83162),
    .in0(net_83115),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79210),
    .ltout(),
    .sr(net_83163)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83162),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_83130),
    .lcout(net_79212),
    .ltout(),
    .sr(net_83163)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83162),
    .in0(gnd),
    .in1(net_83134),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79213),
    .ltout(),
    .sr(net_83163)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83162),
    .in0(net_83157),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79217),
    .ltout(),
    .sr(net_83163)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83285),
    .in0(net_83238),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79333),
    .ltout(),
    .sr(net_83286)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83285),
    .in0(net_83244),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79334),
    .ltout(),
    .sr(net_83286)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83285),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83252_cascademuxed),
    .in3(gnd),
    .lcout(net_79335),
    .ltout(),
    .sr(net_83286)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83285),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83270_cascademuxed),
    .in3(gnd),
    .lcout(net_79338),
    .ltout(),
    .sr(net_83286)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83285),
    .in0(net_83280),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79340),
    .ltout(),
    .sr(net_83286)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83408),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_83376),
    .lcout(net_79458),
    .ltout(),
    .sr(net_83409)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83408),
    .in0(net_83385),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79460),
    .ltout(),
    .sr(net_83409)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83408),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83399_cascademuxed),
    .in3(gnd),
    .lcout(net_79462),
    .ltout(),
    .sr(net_83409)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83531),
    .in0(gnd),
    .in1(net_83509),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79583),
    .ltout(),
    .sr(net_83532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83531),
    .in0(net_83514),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79584),
    .ltout(),
    .sr(net_83532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83531),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83522_cascademuxed),
    .in3(gnd),
    .lcout(net_79585),
    .ltout(),
    .sr(net_83532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83531),
    .in0(net_83526),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79586),
    .ltout(),
    .sr(net_83532)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83654),
    .in0(gnd),
    .in1(net_83614),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79703),
    .ltout(),
    .sr(net_83655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83654),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_83622),
    .lcout(net_79704),
    .ltout(),
    .sr(net_83655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83654),
    .in0(gnd),
    .in1(gnd),
    .in2(net_83627_cascademuxed),
    .in3(gnd),
    .lcout(net_79705),
    .ltout(),
    .sr(net_83655)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83654),
    .in0(net_83649),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79709),
    .ltout(),
    .sr(net_83655)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_8_0 (
    .carryin(t1083),
    .carryout(net_83729),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_83731),
    .in2(net_83732_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_1 (
    .carryin(net_83729),
    .carryout(net_83735),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83737),
    .in2(net_83738_cascademuxed),
    .in3(net_83739),
    .lcout(net_79826),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_2 (
    .carryin(net_83735),
    .carryout(net_83741),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83743),
    .in2(net_83744_cascademuxed),
    .in3(net_83745),
    .lcout(net_79827),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_3 (
    .carryin(net_83741),
    .carryout(net_83747),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83749),
    .in2(net_83750_cascademuxed),
    .in3(net_83751),
    .lcout(net_79828),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_4 (
    .carryin(net_83747),
    .carryout(net_83753),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83755),
    .in2(net_83756_cascademuxed),
    .in3(net_83757),
    .lcout(net_79829),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_5 (
    .carryin(net_83753),
    .carryout(net_83759),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83761),
    .in2(net_83762_cascademuxed),
    .in3(net_83763),
    .lcout(net_79830),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_6 (
    .carryin(net_83759),
    .carryout(net_83765),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83767),
    .in2(net_83768_cascademuxed),
    .in3(net_83769),
    .lcout(net_79831),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_8_7 (
    .carryin(net_83765),
    .carryout(net_83771),
    .ce(),
    .clk(net_83777),
    .in0(gnd),
    .in1(net_83773),
    .in2(net_83774_cascademuxed),
    .in3(net_83775),
    .lcout(net_79832),
    .ltout(),
    .sr(net_83778)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_0 (
    .carryin(net_83815),
    .carryout(net_83852),
    .ce(),
    .clk(net_83900),
    .in0(gnd),
    .in1(net_83854),
    .in2(net_83855_cascademuxed),
    .in3(net_83856),
    .lcout(net_79948),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_1 (
    .carryin(net_83852),
    .carryout(net_83858),
    .ce(),
    .clk(net_83900),
    .in0(gnd),
    .in1(net_83860),
    .in2(net_83861_cascademuxed),
    .in3(net_83862),
    .lcout(net_79949),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_2 (
    .carryin(net_83858),
    .carryout(net_83864),
    .ce(),
    .clk(net_83900),
    .in0(gnd),
    .in1(net_83866),
    .in2(net_83867_cascademuxed),
    .in3(net_83868),
    .lcout(net_79950),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_9_3 (
    .carryin(net_83864),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_83874),
    .lcout(net_79951),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83900),
    .in0(net_83877),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79952),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83900),
    .in0(net_83889),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79954),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_83900),
    .in0(net_83895),
    .in1(gnd),
    .in2(net_83897_cascademuxed),
    .in3(gnd),
    .lcout(net_79955),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_22_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83902),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_86993),
    .in0(gnd),
    .in1(gnd),
    .in2(net_86948_cascademuxed),
    .in3(gnd),
    .lcout(net_83041),
    .ltout(),
    .sr(net_86994)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_86993),
    .in0(gnd),
    .in1(gnd),
    .in2(net_86960_cascademuxed),
    .in3(gnd),
    .lcout(net_83043),
    .ltout(),
    .sr(net_86994)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_86993),
    .in0(gnd),
    .in1(gnd),
    .in2(net_86972_cascademuxed),
    .in3(gnd),
    .lcout(net_83045),
    .ltout(),
    .sr(net_86994)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87116),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87083_cascademuxed),
    .in3(gnd),
    .lcout(net_83166),
    .ltout(),
    .sr(net_87117)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_22_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87116),
    .in0(net_87105),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83170),
    .ltout(),
    .sr(net_87117)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87116),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87113_cascademuxed),
    .in3(gnd),
    .lcout(net_83171),
    .ltout(),
    .sr(net_87117)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_22_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87239),
    .in0(net_87192),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83287),
    .ltout(),
    .sr(net_87240)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_22_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87239),
    .in0(net_87210),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83290),
    .ltout(),
    .sr(net_87240)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87239),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87218_cascademuxed),
    .in3(gnd),
    .lcout(net_83291),
    .ltout(),
    .sr(net_87240)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87239),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87231),
    .lcout(net_83293),
    .ltout(),
    .sr(net_87240)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87239),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87236_cascademuxed),
    .in3(gnd),
    .lcout(net_83294),
    .ltout(),
    .sr(net_87240)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87362),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87342),
    .lcout(net_83414),
    .ltout(),
    .sr(net_87363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87362),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87354),
    .lcout(net_83416),
    .ltout(),
    .sr(net_87363)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87485),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87453),
    .lcout(net_83535),
    .ltout(),
    .sr(net_87486)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87485),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87465),
    .lcout(net_83537),
    .ltout(),
    .sr(net_87486)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_22_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87485),
    .in0(gnd),
    .in1(net_87469),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83538),
    .ltout(),
    .sr(net_87486)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87485),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87483),
    .lcout(net_83540),
    .ltout(),
    .sr(net_87486)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87563_cascademuxed),
    .in3(gnd),
    .lcout(net_83656),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87575_cascademuxed),
    .in3(gnd),
    .lcout(net_83658),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87582),
    .lcout(net_83659),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87588),
    .lcout(net_83660),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87594),
    .lcout(net_83661),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87608),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_87600),
    .lcout(net_83662),
    .ltout(),
    .sr(net_87609)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87731),
    .in0(net_87684),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83779),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87731),
    .in0(net_87702),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83782),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87731),
    .in0(gnd),
    .in1(net_87709),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83783),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87731),
    .in0(gnd),
    .in1(net_87721),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83785),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_87731),
    .in0(gnd),
    .in1(net_87727),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_83786),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_23_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91070),
    .in0(net_91023),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87118),
    .ltout(),
    .sr(net_91071)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_23_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91070),
    .in0(gnd),
    .in1(gnd),
    .in2(net_91031_cascademuxed),
    .in3(gnd),
    .lcout(net_87119),
    .ltout(),
    .sr(net_91071)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_23_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91070),
    .in0(gnd),
    .in1(net_91048),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87122),
    .ltout(),
    .sr(net_91071)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_23_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91070),
    .in0(net_91053),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87123),
    .ltout(),
    .sr(net_91071)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_23_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91070),
    .in0(gnd),
    .in1(gnd),
    .in2(net_91067_cascademuxed),
    .in3(gnd),
    .lcout(net_87125),
    .ltout(),
    .sr(net_91071)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_23_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91193),
    .in0(net_91152),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87242),
    .ltout(),
    .sr(net_91194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_23_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91193),
    .in0(gnd),
    .in1(net_91165),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87244),
    .ltout(),
    .sr(net_91194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_23_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91193),
    .in0(net_91188),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87248),
    .ltout(),
    .sr(net_91194)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_23_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91439),
    .in0(net_91434),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_87494),
    .ltout(),
    .sr(net_91440)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_23_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_91562),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_91536),
    .lcout(net_87613),
    .ltout(),
    .sr(net_91563)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_2_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12452),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8037),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_2_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12464),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8039),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_2_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12475),
    .in1(net_12476),
    .in2(net_12477_cascademuxed),
    .in3(gnd),
    .lcout(net_8041),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12497),
    .clk(net_12498),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12483_cascademuxed),
    .in3(gnd),
    .lcout(net_8042),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_2_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12488),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8043),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12496),
    .lcout(net_8044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_11_0 (
    .carryin(t36),
    .carryout(net_12573),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12575),
    .in2(net_12576_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_1 (
    .carryin(net_12573),
    .carryout(net_12579),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12581),
    .in2(net_12582_cascademuxed),
    .in3(net_12583),
    .lcout(net_8185),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_2 (
    .carryin(net_12579),
    .carryout(net_12585),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12587),
    .in2(net_12588_cascademuxed),
    .in3(net_12589),
    .lcout(net_8186),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_3 (
    .carryin(net_12585),
    .carryout(net_12591),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12593),
    .in2(net_12594_cascademuxed),
    .in3(net_12595),
    .lcout(net_8187),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_4 (
    .carryin(net_12591),
    .carryout(net_12597),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12599),
    .in2(net_12600_cascademuxed),
    .in3(net_12601),
    .lcout(net_8188),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_5 (
    .carryin(net_12597),
    .carryout(net_12603),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12605),
    .in2(net_12606_cascademuxed),
    .in3(net_12607),
    .lcout(net_8189),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_6 (
    .carryin(net_12603),
    .carryout(net_12609),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12611),
    .in2(net_12612_cascademuxed),
    .in3(net_12613),
    .lcout(net_8190),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_11_7 (
    .carryin(net_12609),
    .carryout(net_12615),
    .ce(),
    .clk(net_12621),
    .in0(gnd),
    .in1(net_12617),
    .in2(net_12618_cascademuxed),
    .in3(net_12619),
    .lcout(net_8191),
    .ltout(),
    .sr(net_12622)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_0 (
    .carryin(net_12659),
    .carryout(net_12696),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12698),
    .in2(net_12699_cascademuxed),
    .in3(net_12700),
    .lcout(net_8331),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_1 (
    .carryin(net_12696),
    .carryout(net_12702),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12704),
    .in2(net_12705_cascademuxed),
    .in3(net_12706),
    .lcout(net_8332),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_2 (
    .carryin(net_12702),
    .carryout(net_12708),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12710),
    .in2(net_12711_cascademuxed),
    .in3(net_12712),
    .lcout(net_8333),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_3 (
    .carryin(net_12708),
    .carryout(net_12714),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12716),
    .in2(net_12717_cascademuxed),
    .in3(net_12718),
    .lcout(net_8334),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_4 (
    .carryin(net_12714),
    .carryout(net_12720),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12722),
    .in2(net_12723_cascademuxed),
    .in3(net_12724),
    .lcout(net_8335),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_5 (
    .carryin(net_12720),
    .carryout(net_12726),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12728),
    .in2(net_12729_cascademuxed),
    .in3(net_12730),
    .lcout(net_8336),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_6 (
    .carryin(net_12726),
    .carryout(net_12732),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12734),
    .in2(net_12735_cascademuxed),
    .in3(net_12736),
    .lcout(net_8337),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_12_7 (
    .carryin(net_12732),
    .carryout(net_12738),
    .ce(),
    .clk(net_12744),
    .in0(gnd),
    .in1(net_12740),
    .in2(net_12741_cascademuxed),
    .in3(net_12742),
    .lcout(net_8338),
    .ltout(),
    .sr(net_12745)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(net_12820),
    .in1(gnd),
    .in2(net_12822_cascademuxed),
    .in3(net_12823),
    .lcout(net_8478),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12828_cascademuxed),
    .in3(gnd),
    .lcout(net_8479),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(net_12832),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8480),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12840_cascademuxed),
    .in3(gnd),
    .lcout(net_8481),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(net_12844),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8482),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12853),
    .lcout(net_8483),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(gnd),
    .in1(net_12857),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8484),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12867),
    .in0(gnd),
    .in1(net_12863),
    .in2(gnd),
    .in3(net_12865),
    .lcout(net_8485),
    .ltout(),
    .sr(net_12868)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_14_0 (
    .carryin(t41),
    .carryout(net_12942),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12944),
    .in2(net_12945_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_1 (
    .carryin(net_12942),
    .carryout(net_12948),
    .ce(),
    .clk(net_12990),
    .in0(gnd),
    .in1(net_12950),
    .in2(net_12951_cascademuxed),
    .in3(net_12952),
    .lcout(net_8626),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(gnd),
    .in1(net_12956),
    .in2(net_12957_cascademuxed),
    .in3(net_12958),
    .lcout(net_8627),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(gnd),
    .in1(net_12962),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8628),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(net_12967),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8629),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12975_cascademuxed),
    .in3(gnd),
    .lcout(net_8630),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(net_12979),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12982),
    .lcout(net_8631),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12990),
    .in0(net_12985),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8632),
    .ltout(),
    .sr(net_12991)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_15_0 (
    .carryin(t46),
    .carryout(net_13065),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_13067),
    .in2(net_13068_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_2_15_1 (
    .carryin(net_13065),
    .carryout(net_13071),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_13073),
    .in2(net_13074_cascademuxed),
    .in3(net_13075),
    .lcout(net_8773),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001011001101001),
    .SEQ_MODE(4'b0000)
  ) lc40_2_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_13079),
    .in2(net_13080_cascademuxed),
    .in3(net_13081),
    .lcout(net_8774),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_2_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_13084),
    .in1(net_13085),
    .in2(net_13086_cascademuxed),
    .in3(gnd),
    .lcout(net_8775),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13113),
    .in0(net_13090),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8776),
    .ltout(),
    .sr(net_13114)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13113),
    .in0(gnd),
    .in1(net_13097),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8777),
    .ltout(),
    .sr(net_13114)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13113),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13105),
    .lcout(net_8778),
    .ltout(),
    .sr(net_13114)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13113),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13111),
    .lcout(net_8779),
    .ltout(),
    .sr(net_13114)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13236),
    .in0(net_13189),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8919),
    .ltout(),
    .sr(net_13237)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13236),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13198),
    .lcout(net_8920),
    .ltout(),
    .sr(net_13237)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13236),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13203_cascademuxed),
    .in3(gnd),
    .lcout(net_8921),
    .ltout(),
    .sr(net_13237)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13236),
    .in0(net_13207),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8922),
    .ltout(),
    .sr(net_13237)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_2_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_13214),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8923),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_2_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_13219),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_8924),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13227_cascademuxed),
    .in3(gnd),
    .lcout(net_8925),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13233_cascademuxed),
    .in3(gnd),
    .lcout(net_8926),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13359),
    .in0(net_13324),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9068),
    .ltout(),
    .sr(net_13360)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13359),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13345),
    .lcout(net_9071),
    .ltout(),
    .sr(net_13360)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13359),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13356_cascademuxed),
    .in3(gnd),
    .lcout(net_9073),
    .ltout(),
    .sr(net_13360)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13482),
    .in0(gnd),
    .in1(net_13436),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9213),
    .ltout(),
    .sr(net_13483)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13482),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13444),
    .lcout(net_9214),
    .ltout(),
    .sr(net_13483)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13482),
    .in0(gnd),
    .in1(net_13460),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9217),
    .ltout(),
    .sr(net_13483)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13482),
    .in0(gnd),
    .in1(net_13472),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9219),
    .ltout(),
    .sr(net_13483)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13482),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13479_cascademuxed),
    .in3(gnd),
    .lcout(net_9220),
    .ltout(),
    .sr(net_13483)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13560_cascademuxed),
    .in3(gnd),
    .lcout(net_9360),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13567),
    .lcout(net_9361),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(net_13576),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9363),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(gnd),
    .in1(net_13583),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9364),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13591),
    .lcout(net_9365),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13596_cascademuxed),
    .in3(gnd),
    .lcout(net_9366),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13605),
    .in0(net_13600),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9367),
    .ltout(),
    .sr(net_13606)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010001001110111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_1_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11304),
    .in1(net_11305),
    .in2(gnd),
    .in3(net_11307),
    .lcout(net_6673),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_1_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11351),
    .in0(net_11310),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_6674),
    .ltout(),
    .sr(net_11352)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11322),
    .in1(net_11323),
    .in2(net_11324_cascademuxed),
    .in3(net_11325),
    .lcout(net_6676),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11336_cascademuxed),
    .in3(gnd),
    .lcout(net_6678),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010010110100101),
    .SEQ_MODE(4'b0000)
  ) lc40_2_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11346),
    .in1(gnd),
    .in2(net_11348_cascademuxed),
    .in3(gnd),
    .lcout(net_6680),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13728),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13690),
    .lcout(net_9508),
    .ltout(),
    .sr(net_13729)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_20_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13728),
    .in0(gnd),
    .in1(net_13700),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9510),
    .ltout(),
    .sr(net_13729)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_20_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13728),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_13708),
    .lcout(net_9511),
    .ltout(),
    .sr(net_13729)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13728),
    .in0(net_13711),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9512),
    .ltout(),
    .sr(net_13729)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13728),
    .in0(net_13723),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9514),
    .ltout(),
    .sr(net_13729)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_21_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13851),
    .in0(net_13810),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9655),
    .ltout(),
    .sr(net_13852)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_21_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13851),
    .in0(gnd),
    .in1(net_13829),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9658),
    .ltout(),
    .sr(net_13852)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_22_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13974),
    .in0(gnd),
    .in1(net_13928),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9801),
    .ltout(),
    .sr(net_13975)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_22_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_13974),
    .in0(gnd),
    .in1(gnd),
    .in2(net_13959_cascademuxed),
    .in3(gnd),
    .lcout(net_9806),
    .ltout(),
    .sr(net_13975)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_23_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_14097),
    .in0(net_14074),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_9952),
    .ltout(),
    .sr(net_14098)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11514),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11469_cascademuxed),
    .in3(gnd),
    .lcout(net_6825),
    .ltout(),
    .sr(net_11515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000110000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_11474),
    .in2(net_11475_cascademuxed),
    .in3(net_11476),
    .lcout(net_6826),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000110000100),
    .SEQ_MODE(4'b0000)
  ) lc40_2_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11479),
    .in1(net_11480),
    .in2(net_11481_cascademuxed),
    .in3(net_11482),
    .lcout(net_6827),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11514),
    .in0(net_11485),
    .in1(net_11486),
    .in2(net_11487_cascademuxed),
    .in3(net_11488),
    .lcout(net_6828),
    .ltout(),
    .sr(net_11515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11514),
    .in0(gnd),
    .in1(net_11492),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_6829),
    .ltout(),
    .sr(net_11515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001000000001001),
    .SEQ_MODE(4'b0000)
  ) lc40_2_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11497),
    .in1(net_11498),
    .in2(net_11499_cascademuxed),
    .in3(net_11500),
    .lcout(net_6830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11503),
    .in1(gnd),
    .in2(net_11505_cascademuxed),
    .in3(net_11506),
    .lcout(net_6831),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100010111000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11509),
    .in1(net_11510),
    .in2(net_11511_cascademuxed),
    .in3(gnd),
    .lcout(net_6832),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100000100010),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11590),
    .in1(net_11591),
    .in2(gnd),
    .in3(net_11593),
    .lcout(net_7008),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000010000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11596),
    .in1(net_11597),
    .in2(net_11598_cascademuxed),
    .in3(gnd),
    .lcout(net_7009),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11637),
    .in0(gnd),
    .in1(net_11603),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7010),
    .ltout(),
    .sr(net_11638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11637),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_11611),
    .lcout(net_7011),
    .ltout(),
    .sr(net_11638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010010000100),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11614),
    .in1(net_11615),
    .in2(net_11616_cascademuxed),
    .in3(gnd),
    .lcout(net_7012),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010001011110011),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11620),
    .in1(net_11621),
    .in2(net_11622_cascademuxed),
    .in3(net_11623),
    .lcout(net_7013),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11626),
    .in1(net_11627),
    .in2(net_11628_cascademuxed),
    .in3(net_11629),
    .lcout(net_7014),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111101000101),
    .SEQ_MODE(4'b0000)
  ) lc40_2_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11632),
    .in1(net_11633),
    .in2(net_11634_cascademuxed),
    .in3(net_11635),
    .lcout(net_7015),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11713),
    .in1(net_11714),
    .in2(net_11715_cascademuxed),
    .in3(net_11716),
    .lcout(net_7155),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111001000100),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11719),
    .in1(net_11720),
    .in2(gnd),
    .in3(net_11722),
    .lcout(net_7156),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_11728),
    .lcout(net_7157),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001000000001001),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11731),
    .in1(net_11732),
    .in2(net_11733_cascademuxed),
    .in3(net_11734),
    .lcout(net_7158),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000100001),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11737),
    .in1(net_11738),
    .in2(net_11739_cascademuxed),
    .in3(net_11740),
    .lcout(net_7159),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11760),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11745_cascademuxed),
    .in3(gnd),
    .lcout(net_7160),
    .ltout(),
    .sr(net_11761)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011100010),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11749),
    .in1(net_11750),
    .in2(net_11751_cascademuxed),
    .in3(gnd),
    .lcout(net_7161),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11755),
    .in1(net_11756),
    .in2(gnd),
    .in3(net_11758),
    .lcout(net_7162),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11883),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11838_cascademuxed),
    .in3(gnd),
    .lcout(net_7302),
    .ltout(),
    .sr(net_11884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_11848),
    .in1(gnd),
    .in2(net_11850_cascademuxed),
    .in3(net_11851),
    .lcout(net_7304),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11883),
    .in0(gnd),
    .in1(net_11855),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7305),
    .ltout(),
    .sr(net_11884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11883),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11862_cascademuxed),
    .in3(gnd),
    .lcout(net_7306),
    .ltout(),
    .sr(net_11884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11883),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_11875),
    .lcout(net_7308),
    .ltout(),
    .sr(net_11884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_11883),
    .in0(net_11878),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7309),
    .ltout(),
    .sr(net_11884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_11962),
    .lcout(net_7449),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11967_cascademuxed),
    .in3(gnd),
    .lcout(net_7450),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11973_cascademuxed),
    .in3(gnd),
    .lcout(net_7451),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11979_cascademuxed),
    .in3(gnd),
    .lcout(net_7452),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(net_11983),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7453),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(gnd),
    .in1(gnd),
    .in2(net_11991_cascademuxed),
    .in3(gnd),
    .lcout(net_7454),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12006),
    .in0(net_11995),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7455),
    .ltout(),
    .sr(net_12007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_2_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12128),
    .clk(net_12129),
    .in0(gnd),
    .in1(net_12083),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7596),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_2_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12088),
    .in1(net_12089),
    .in2(net_12090_cascademuxed),
    .in3(net_12091),
    .lcout(net_7597),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12128),
    .clk(net_12129),
    .in0(net_12100),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7599),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12128),
    .clk(net_12129),
    .in0(net_12106),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7600),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12128),
    .clk(net_12129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12120_cascademuxed),
    .in3(gnd),
    .lcout(net_7602),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12128),
    .clk(net_12129),
    .in0(net_12124),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7603),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12205),
    .in1(net_12206),
    .in2(net_12207_cascademuxed),
    .in3(net_12208),
    .lcout(net_7743),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12211),
    .in1(net_12212),
    .in2(net_12213_cascademuxed),
    .in3(net_12214),
    .lcout(net_7744),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12251),
    .clk(net_12252),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12220),
    .lcout(net_7745),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101011010000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12223),
    .in1(net_12224),
    .in2(net_12225_cascademuxed),
    .in3(net_12226),
    .lcout(net_7746),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12229),
    .in1(net_12230),
    .in2(net_12231_cascademuxed),
    .in3(net_12232),
    .lcout(net_7747),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12251),
    .clk(net_12252),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12238),
    .lcout(net_7748),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12251),
    .clk(net_12252),
    .in0(net_12241),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7749),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_12251),
    .clk(net_12252),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12249_cascademuxed),
    .in3(gnd),
    .lcout(net_7750),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(net_12328),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7890),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_2_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12334),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7891),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12343),
    .lcout(net_7892),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(net_12346),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7893),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(net_12352),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7894),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(net_12358),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7895),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(net_12364),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_7896),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_2_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12375),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_12373),
    .lcout(net_7897),
    .ltout(),
    .sr(net_12376)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(net_16283),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12377),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16291),
    .lcout(net_12378),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16296_cascademuxed),
    .in3(gnd),
    .lcout(net_12379),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(net_16300),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12380),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16309),
    .lcout(net_12381),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16315),
    .lcout(net_12382),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16320_cascademuxed),
    .in3(gnd),
    .lcout(net_12383),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16329),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16326_cascademuxed),
    .in3(gnd),
    .lcout(net_12384),
    .ltout(),
    .sr(net_16330)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(net_16406),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12500),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16414),
    .lcout(net_12501),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16419_cascademuxed),
    .in3(gnd),
    .lcout(net_12502),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16425_cascademuxed),
    .in3(gnd),
    .lcout(net_12503),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16431_cascademuxed),
    .in3(gnd),
    .lcout(net_12504),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(net_16436),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12505),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16452),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16443_cascademuxed),
    .in3(gnd),
    .lcout(net_12506),
    .ltout(),
    .sr(net_16453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16450),
    .lcout(net_12507),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_0 (
    .carryin(t106),
    .carryout(net_16527),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16529),
    .in2(net_16530_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_1 (
    .carryin(net_16527),
    .carryout(net_16533),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16535),
    .in2(net_16536_cascademuxed),
    .in3(net_16537),
    .lcout(net_12624),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_2 (
    .carryin(net_16533),
    .carryout(net_16539),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16541),
    .in2(net_16542_cascademuxed),
    .in3(net_16543),
    .lcout(net_12625),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_3 (
    .carryin(net_16539),
    .carryout(net_16545),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16547),
    .in2(net_16548_cascademuxed),
    .in3(net_16549),
    .lcout(net_12626),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_4 (
    .carryin(net_16545),
    .carryout(net_16551),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16553),
    .in2(net_16554_cascademuxed),
    .in3(net_16555),
    .lcout(net_12627),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_5 (
    .carryin(net_16551),
    .carryout(net_16557),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16559),
    .in2(net_16560_cascademuxed),
    .in3(net_16561),
    .lcout(net_12628),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_6 (
    .carryin(net_16557),
    .carryout(net_16563),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16565),
    .in2(net_16566_cascademuxed),
    .in3(net_16567),
    .lcout(net_12629),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16573),
    .lcout(net_12630),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_13_0 (
    .carryin(t116),
    .carryout(net_16650),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16652),
    .in2(net_16653_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_1 (
    .carryin(net_16650),
    .carryout(net_16656),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16658),
    .in2(net_16659_cascademuxed),
    .in3(net_16660),
    .lcout(net_12747),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_2 (
    .carryin(net_16656),
    .carryout(net_16662),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16664),
    .in2(net_16665_cascademuxed),
    .in3(net_16666),
    .lcout(net_12748),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_3 (
    .carryin(net_16662),
    .carryout(net_16668),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16670),
    .in2(net_16671_cascademuxed),
    .in3(net_16672),
    .lcout(net_12749),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_4 (
    .carryin(net_16668),
    .carryout(net_16674),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16676),
    .in2(net_16677_cascademuxed),
    .in3(net_16678),
    .lcout(net_12750),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_5 (
    .carryin(net_16674),
    .carryout(net_16680),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16682),
    .in2(net_16683_cascademuxed),
    .in3(net_16684),
    .lcout(net_12751),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_6 (
    .carryin(net_16680),
    .carryout(net_16686),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16688),
    .in2(net_16689_cascademuxed),
    .in3(net_16690),
    .lcout(net_12752),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_7 (
    .carryin(net_16686),
    .carryout(net_16692),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16694),
    .in2(net_16695_cascademuxed),
    .in3(net_16696),
    .lcout(net_12753),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_0 (
    .carryin(net_16736),
    .carryout(net_16773),
    .ce(),
    .clk(net_16821),
    .in0(gnd),
    .in1(net_16775),
    .in2(net_16776_cascademuxed),
    .in3(net_16777),
    .lcout(net_12869),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16821),
    .in0(net_16780),
    .in1(gnd),
    .in2(net_16782_cascademuxed),
    .in3(net_16783),
    .lcout(net_12870),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16821),
    .in0(gnd),
    .in1(net_16787),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12871),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16794_cascademuxed),
    .in3(gnd),
    .lcout(net_12872),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16821),
    .in0(gnd),
    .in1(net_16799),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12873),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_16804),
    .in1(net_16805),
    .in2(gnd),
    .in3(net_16807),
    .lcout(net_12874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16821),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16812_cascademuxed),
    .in3(gnd),
    .lcout(net_12875),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16821),
    .in0(gnd),
    .in1(net_16817),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12876),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_0 (
    .carryin(t126),
    .carryout(net_16896),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16898),
    .in2(net_16899_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_1 (
    .carryin(net_16896),
    .carryout(net_16902),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16904),
    .in2(net_16905_cascademuxed),
    .in3(net_16906),
    .lcout(net_12993),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_2 (
    .carryin(net_16902),
    .carryout(net_16908),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16910),
    .in2(net_16911_cascademuxed),
    .in3(net_16912),
    .lcout(net_12994),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_3 (
    .carryin(net_16908),
    .carryout(net_16914),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16916),
    .in2(net_16917_cascademuxed),
    .in3(net_16918),
    .lcout(net_12995),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_4 (
    .carryin(net_16914),
    .carryout(net_16920),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16922),
    .in2(net_16923_cascademuxed),
    .in3(net_16924),
    .lcout(net_12996),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_5 (
    .carryin(net_16920),
    .carryout(net_16926),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16928),
    .in2(net_16929_cascademuxed),
    .in3(net_16930),
    .lcout(net_12997),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_6 (
    .carryin(net_16926),
    .carryout(net_16932),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16934),
    .in2(net_16935_cascademuxed),
    .in3(net_16936),
    .lcout(net_12998),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16942),
    .lcout(net_12999),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17023),
    .lcout(net_13115),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17029),
    .lcout(net_13116),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17033),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13117),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17041),
    .lcout(net_13118),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17045),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13119),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17067),
    .in0(gnd),
    .in1(net_17051),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13120),
    .ltout(),
    .sr(net_17068)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_3_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17057),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13121),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17067),
    .in0(net_17062),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13122),
    .ltout(),
    .sr(net_17068)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(net_17143),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13238),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17158),
    .lcout(net_13240),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17164),
    .lcout(net_13241),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17169_cascademuxed),
    .in3(gnd),
    .lcout(net_13242),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(net_17173),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13243),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17190),
    .in0(net_17179),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13244),
    .ltout(),
    .sr(net_17191)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_3_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_17185),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13245),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_17312),
    .clk(net_17313),
    .in0(net_17266),
    .in1(net_17267),
    .in2(net_17268_cascademuxed),
    .in3(net_17269),
    .lcout(net_13361),
    .ltout(),
    .sr(net_17314)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_3_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17291),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13365),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_17312),
    .clk(net_17313),
    .in0(net_17296),
    .in1(net_17297),
    .in2(net_17298_cascademuxed),
    .in3(net_17299),
    .lcout(net_13366),
    .ltout(),
    .sr(net_17314)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_17312),
    .clk(net_17313),
    .in0(net_17302),
    .in1(net_17303),
    .in2(net_17304_cascademuxed),
    .in3(net_17305),
    .lcout(net_13367),
    .ltout(),
    .sr(net_17314)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_3_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17309),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13368),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(net_17402),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13486),
    .ltout(),
    .sr(net_17437)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17421_cascademuxed),
    .in3(gnd),
    .lcout(net_13489),
    .ltout(),
    .sr(net_17437)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_1_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15135),
    .in1(net_15136),
    .in2(net_15137_cascademuxed),
    .in3(net_15138),
    .lcout(net_11229),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110011101100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_1_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15181),
    .clk(net_15182),
    .in0(net_15141),
    .in1(net_15142),
    .in2(net_15143_cascademuxed),
    .in3(gnd),
    .lcout(net_11230),
    .ltout(),
    .sr(net_15183)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_1_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15181),
    .clk(net_15182),
    .in0(net_15147),
    .in1(net_15148),
    .in2(net_15149_cascademuxed),
    .in3(net_15150),
    .lcout(net_11231),
    .ltout(),
    .sr(net_15183)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15181),
    .clk(net_15182),
    .in0(net_15153),
    .in1(net_15154),
    .in2(net_15155_cascademuxed),
    .in3(net_15156),
    .lcout(net_11232),
    .ltout(),
    .sr(net_15183)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000101000001010),
    .SEQ_MODE(4'b0000)
  ) lc40_3_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15171),
    .in1(gnd),
    .in2(net_15173_cascademuxed),
    .in3(gnd),
    .lcout(net_11235),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010111000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15181),
    .clk(net_15182),
    .in0(net_15177),
    .in1(net_15178),
    .in2(net_15179_cascademuxed),
    .in3(net_15180),
    .lcout(net_11236),
    .ltout(),
    .sr(net_15183)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_17521),
    .lcout(net_13608),
    .ltout(),
    .sr(net_17560)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_21_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17682),
    .in0(gnd),
    .in1(net_17666),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13735),
    .ltout(),
    .sr(net_17683)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_21_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17682),
    .in0(net_17671),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13736),
    .ltout(),
    .sr(net_17683)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_22_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17805),
    .in0(gnd),
    .in1(net_17777),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_13856),
    .ltout(),
    .sr(net_17806)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100101000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15298),
    .in1(net_15299),
    .in2(net_15300_cascademuxed),
    .in3(net_15301),
    .lcout(net_11357),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000010100000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15304),
    .in1(net_15305),
    .in2(net_15306_cascademuxed),
    .in3(net_15307),
    .lcout(net_11358),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15344),
    .clk(net_15345),
    .in0(gnd),
    .in1(net_15311),
    .in2(net_15312_cascademuxed),
    .in3(net_15313),
    .lcout(net_11359),
    .ltout(),
    .sr(net_15346)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100011000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15316),
    .in1(net_15317),
    .in2(net_15318_cascademuxed),
    .in3(net_15319),
    .lcout(net_11360),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15344),
    .clk(net_15345),
    .in0(net_15322),
    .in1(net_15323),
    .in2(gnd),
    .in3(net_15325),
    .lcout(net_11361),
    .ltout(),
    .sr(net_15346)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010001010000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15328),
    .in1(net_15329),
    .in2(net_15330_cascademuxed),
    .in3(net_15331),
    .lcout(net_11362),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111001100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15344),
    .clk(net_15345),
    .in0(gnd),
    .in1(net_15335),
    .in2(gnd),
    .in3(net_15337),
    .lcout(net_11363),
    .ltout(),
    .sr(net_15346)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110011001100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15344),
    .clk(net_15345),
    .in0(gnd),
    .in1(net_15341),
    .in2(net_15342_cascademuxed),
    .in3(net_15343),
    .lcout(net_11364),
    .ltout(),
    .sr(net_15346)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100011000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15421),
    .in1(net_15422),
    .in2(net_15423_cascademuxed),
    .in3(net_15424),
    .lcout(net_11516),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15427),
    .in1(net_15428),
    .in2(net_15429_cascademuxed),
    .in3(net_15430),
    .lcout(net_11517),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111011101110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15467),
    .clk(net_15468),
    .in0(net_15433),
    .in1(net_15434),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11518),
    .ltout(),
    .sr(net_15469)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000111110001000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15467),
    .clk(net_15468),
    .in0(net_15439),
    .in1(net_15440),
    .in2(net_15441_cascademuxed),
    .in3(net_15442),
    .lcout(net_11519),
    .ltout(),
    .sr(net_15469)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110100000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15467),
    .clk(net_15468),
    .in0(net_15445),
    .in1(gnd),
    .in2(net_15447_cascademuxed),
    .in3(net_15448),
    .lcout(net_11520),
    .ltout(),
    .sr(net_15469)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010101001111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15451),
    .in1(net_15452),
    .in2(net_15453_cascademuxed),
    .in3(net_15454),
    .lcout(net_11521),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101000010000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15457),
    .in1(net_15458),
    .in2(net_15459_cascademuxed),
    .in3(net_15460),
    .lcout(net_11522),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15463),
    .in1(net_15464),
    .in2(net_15465_cascademuxed),
    .in3(net_15466),
    .lcout(net_11523),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110001000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15591),
    .in0(net_15544),
    .in1(net_15545),
    .in2(net_15546_cascademuxed),
    .in3(net_15547),
    .lcout(net_11639),
    .ltout(),
    .sr(net_15592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111011101110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15556),
    .in1(net_15557),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11641),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15591),
    .in0(gnd),
    .in1(gnd),
    .in2(net_15564_cascademuxed),
    .in3(gnd),
    .lcout(net_11642),
    .ltout(),
    .sr(net_15592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010011100100111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15568),
    .in1(net_15569),
    .in2(net_15570_cascademuxed),
    .in3(gnd),
    .lcout(net_11643),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000100010),
    .SEQ_MODE(4'b0000)
  ) lc40_3_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15574),
    .in1(net_15575),
    .in2(gnd),
    .in3(net_15577),
    .lcout(net_11644),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15591),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_15583),
    .lcout(net_11645),
    .ltout(),
    .sr(net_15592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_15587),
    .in2(gnd),
    .in3(net_15589),
    .lcout(net_11646),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_15668),
    .in2(gnd),
    .in3(net_15670),
    .lcout(net_11762),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(gnd),
    .in1(net_15674),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11763),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_15682),
    .lcout(net_11764),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(gnd),
    .in1(net_15692),
    .in2(gnd),
    .in3(net_15694),
    .lcout(net_11766),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(net_15697),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11767),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(gnd),
    .in1(gnd),
    .in2(net_15705_cascademuxed),
    .in3(gnd),
    .lcout(net_11768),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15714),
    .in0(net_15709),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11769),
    .ltout(),
    .sr(net_15715)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15836),
    .clk(net_15837),
    .in0(gnd),
    .in1(net_15791),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11885),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15836),
    .clk(net_15837),
    .in0(gnd),
    .in1(net_15797),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11886),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15836),
    .clk(net_15837),
    .in0(net_15808),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11888),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101001001010),
    .SEQ_MODE(4'b0000)
  ) lc40_3_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_15814),
    .in1(net_15815),
    .in2(net_15816_cascademuxed),
    .in3(net_15817),
    .lcout(net_11889),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_3_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15836),
    .clk(net_15837),
    .in0(net_15820),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_11890),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_15827),
    .in2(net_15828_cascademuxed),
    .in3(net_15829),
    .lcout(net_11891),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_15836),
    .clk(net_15837),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_15835),
    .lcout(net_11892),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_7_0 (
    .carryin(t85),
    .carryout(net_15912),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_15914),
    .in2(net_15915_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_1 (
    .carryin(net_15912),
    .carryout(net_15918),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15920),
    .in2(net_15921_cascademuxed),
    .in3(net_15922),
    .lcout(net_12009),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_2 (
    .carryin(net_15918),
    .carryout(net_15924),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15926),
    .in2(net_15927_cascademuxed),
    .in3(net_15928),
    .lcout(net_12010),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_3 (
    .carryin(net_15924),
    .carryout(net_15930),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15932),
    .in2(net_15933_cascademuxed),
    .in3(net_15934),
    .lcout(net_12011),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_4 (
    .carryin(net_15930),
    .carryout(net_15936),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15938),
    .in2(net_15939_cascademuxed),
    .in3(net_15940),
    .lcout(net_12012),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_5 (
    .carryin(net_15936),
    .carryout(net_15942),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15944),
    .in2(net_15945_cascademuxed),
    .in3(net_15946),
    .lcout(net_12013),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_7_6 (
    .carryin(net_15942),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_15952),
    .lcout(net_12014),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15960),
    .in0(gnd),
    .in1(net_15956),
    .in2(net_15957_cascademuxed),
    .in3(gnd),
    .lcout(net_12015),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_16082),
    .clk(net_16083),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16038_cascademuxed),
    .in3(gnd),
    .lcout(net_12131),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_3_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_16082),
    .clk(net_16083),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16051),
    .lcout(net_12133),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_16060),
    .in1(net_16061),
    .in2(gnd),
    .in3(net_16063),
    .lcout(net_12135),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_3_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_16082),
    .clk(net_16083),
    .in0(gnd),
    .in1(net_16079),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12138),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_0 (
    .carryin(t94),
    .carryout(net_16158),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16160),
    .in2(net_16161_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_1 (
    .carryin(net_16158),
    .carryout(net_16164),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16166),
    .in2(net_16167_cascademuxed),
    .in3(net_16168),
    .lcout(net_12255),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_2 (
    .carryin(net_16164),
    .carryout(net_16170),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16172),
    .in2(net_16173_cascademuxed),
    .in3(net_16174),
    .lcout(net_12256),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_3 (
    .carryin(net_16170),
    .carryout(net_16176),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16178),
    .in2(net_16179_cascademuxed),
    .in3(net_16180),
    .lcout(net_12257),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_4 (
    .carryin(net_16176),
    .carryout(net_16182),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16184),
    .in2(net_16185_cascademuxed),
    .in3(net_16186),
    .lcout(net_12258),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_5 (
    .carryin(net_16182),
    .carryout(net_16188),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16190),
    .in2(net_16191_cascademuxed),
    .in3(net_16192),
    .lcout(net_12259),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_6 (
    .carryin(net_16188),
    .carryout(net_16194),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16196),
    .in2(net_16197_cascademuxed),
    .in3(net_16198),
    .lcout(net_12260),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_3_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_16204),
    .lcout(net_12261),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_0 (
    .carryin(net_20075),
    .carryout(net_20112),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20114),
    .in2(net_20115_cascademuxed),
    .in3(net_20116),
    .lcout(net_16208),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_1 (
    .carryin(net_20112),
    .carryout(net_20118),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20120),
    .in2(net_20121_cascademuxed),
    .in3(net_20122),
    .lcout(net_16209),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_2 (
    .carryin(net_20118),
    .carryout(net_20124),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20126),
    .in2(net_20127_cascademuxed),
    .in3(net_20128),
    .lcout(net_16210),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_3 (
    .carryin(net_20124),
    .carryout(net_20130),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20132),
    .in2(net_20133_cascademuxed),
    .in3(net_20134),
    .lcout(net_16211),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_4 (
    .carryin(net_20130),
    .carryout(net_20136),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20138),
    .in2(net_20139_cascademuxed),
    .in3(net_20140),
    .lcout(net_16212),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_5 (
    .carryin(net_20136),
    .carryout(net_20142),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20144),
    .in2(net_20145_cascademuxed),
    .in3(net_20146),
    .lcout(net_16213),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_6 (
    .carryin(net_20142),
    .carryout(net_20148),
    .ce(),
    .clk(net_20160),
    .in0(gnd),
    .in1(net_20150),
    .in2(net_20151_cascademuxed),
    .in3(net_20152),
    .lcout(net_16214),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20160),
    .in0(net_20155),
    .in1(net_20156),
    .in2(gnd),
    .in3(net_20158),
    .lcout(net_16215),
    .ltout(),
    .sr(net_20161)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(net_20237),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16331),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(net_20242),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16332),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20251),
    .lcout(net_16333),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(net_20255),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16334),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20262_cascademuxed),
    .in3(gnd),
    .lcout(net_16335),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(net_20266),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16336),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20274_cascademuxed),
    .in3(gnd),
    .lcout(net_16337),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20283),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20281),
    .lcout(net_16338),
    .ltout(),
    .sr(net_20284)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_20405),
    .clk(net_20406),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20362),
    .lcout(net_16454),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_20405),
    .clk(net_20406),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20367_cascademuxed),
    .in3(gnd),
    .lcout(net_16455),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_4_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_20371),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16456),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_20405),
    .clk(net_20406),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20380),
    .lcout(net_16457),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_4_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_20383),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16458),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_20405),
    .clk(net_20406),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20391_cascademuxed),
    .in3(gnd),
    .lcout(net_16459),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_20405),
    .clk(net_20406),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20404),
    .lcout(net_16461),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_0 (
    .carryin(t207),
    .carryout(t209),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20483),
    .in2(net_20484_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_1 (
    .carryin(t209),
    .carryout(t210),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20489),
    .in2(net_20490_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_2 (
    .carryin(t210),
    .carryout(t211),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20495),
    .in2(net_20496_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_3 (
    .carryin(t211),
    .carryout(t212),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20501),
    .in2(net_20502_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_4 (
    .carryin(t212),
    .carryout(t213),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20507),
    .in2(net_20508_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_5 (
    .carryin(t213),
    .carryout(t214),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20513),
    .in2(net_20514_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_6 (
    .carryin(t214),
    .carryout(net_20517),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_20519),
    .in2(net_20520_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_13_7 (
    .carryin(net_20517),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20527),
    .lcout(net_16584),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(gnd),
    .in1(net_20606),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16700),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(net_20611),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16701),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20625_cascademuxed),
    .in3(gnd),
    .lcout(net_16703),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(net_20629),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16704),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20637_cascademuxed),
    .in3(gnd),
    .lcout(net_16705),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20644),
    .lcout(net_16706),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20652),
    .in0(net_20647),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16707),
    .ltout(),
    .sr(net_20653)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(net_20728),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16823),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20737),
    .lcout(net_16824),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20743),
    .lcout(net_16825),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(net_20746),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16826),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(net_20752),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16827),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(gnd),
    .in1(net_20759),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16828),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20766_cascademuxed),
    .in3(gnd),
    .lcout(net_16829),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20775),
    .in0(net_20770),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16830),
    .ltout(),
    .sr(net_20776)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(net_20852),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16946),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(net_20858),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16947),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20877_cascademuxed),
    .in3(gnd),
    .lcout(net_16950),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20883_cascademuxed),
    .in3(gnd),
    .lcout(net_16951),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(net_20888),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_16952),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20898),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20896),
    .lcout(net_16953),
    .ltout(),
    .sr(net_20899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20977),
    .lcout(net_17069),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(net_20980),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_17070),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(net_20993),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_17072),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_21001),
    .lcout(net_17073),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(gnd),
    .in2(net_21006_cascademuxed),
    .in3(gnd),
    .lcout(net_17074),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_21013),
    .lcout(net_17075),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21021),
    .in0(gnd),
    .in1(net_21017),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_17076),
    .ltout(),
    .sr(net_21022)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_21143),
    .clk(net_21144),
    .in0(net_21115),
    .in1(net_21116),
    .in2(net_21117_cascademuxed),
    .in3(net_21118),
    .lcout(net_17195),
    .ltout(),
    .sr(net_21145)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21267),
    .in0(gnd),
    .in1(gnd),
    .in2(net_21222_cascademuxed),
    .in3(gnd),
    .lcout(net_17315),
    .ltout(),
    .sr(net_21268)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21267),
    .in0(gnd),
    .in1(gnd),
    .in2(net_21258_cascademuxed),
    .in3(gnd),
    .lcout(net_17321),
    .ltout(),
    .sr(net_21268)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21267),
    .in0(gnd),
    .in1(gnd),
    .in2(net_21264_cascademuxed),
    .in3(gnd),
    .lcout(net_17322),
    .ltout(),
    .sr(net_21268)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010111110101),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_18966),
    .in1(net_18967),
    .in2(net_18968_cascademuxed),
    .in3(net_18969),
    .lcout(net_15060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101011111010),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_18978),
    .in1(gnd),
    .in2(net_18980_cascademuxed),
    .in3(gnd),
    .lcout(net_15062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_18984),
    .in1(net_18985),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15063),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011101010),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_18990),
    .in1(net_18991),
    .in2(net_18992_cascademuxed),
    .in3(net_18993),
    .lcout(net_15064),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111010101010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19012),
    .clk(net_19013),
    .in0(net_18996),
    .in1(net_18997),
    .in2(net_18998_cascademuxed),
    .in3(net_18999),
    .lcout(net_15065),
    .ltout(),
    .sr(net_19014)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010101001111111),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19002),
    .in1(net_19003),
    .in2(net_19004_cascademuxed),
    .in3(net_19005),
    .lcout(net_15066),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100011111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_4_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19008),
    .in1(net_19009),
    .in2(net_19010_cascademuxed),
    .in3(net_19011),
    .lcout(net_15067),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_20_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21390),
    .in0(gnd),
    .in1(net_21368),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_17442),
    .ltout(),
    .sr(net_21391)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21390),
    .in0(gnd),
    .in1(gnd),
    .in2(net_21375_cascademuxed),
    .in3(gnd),
    .lcout(net_17443),
    .ltout(),
    .sr(net_21391)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_22_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21636),
    .in0(gnd),
    .in1(net_21626),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_17690),
    .ltout(),
    .sr(net_21637)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_0 (
    .carryin(t146),
    .carryout(net_19128),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19130),
    .in2(net_19131_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_1 (
    .carryin(net_19128),
    .carryout(net_19134),
    .ce(),
    .clk(gnd),
    .in0(net_19135),
    .in1(net_19136),
    .in2(net_19137_cascademuxed),
    .in3(net_19138),
    .lcout(net_15189),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_2 (
    .carryin(net_19134),
    .carryout(net_19140),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19142),
    .in2(net_19143_cascademuxed),
    .in3(net_19144),
    .lcout(net_15190),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_3 (
    .carryin(net_19140),
    .carryout(net_19146),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19148),
    .in2(net_19149_cascademuxed),
    .in3(net_19150),
    .lcout(net_15191),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_4 (
    .carryin(net_19146),
    .carryout(net_19152),
    .ce(),
    .clk(gnd),
    .in0(net_19153),
    .in1(net_19154),
    .in2(net_19155_cascademuxed),
    .in3(net_19156),
    .lcout(net_15192),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_5 (
    .carryin(net_19152),
    .carryout(net_19158),
    .ce(),
    .clk(gnd),
    .in0(net_19159),
    .in1(net_19160),
    .in2(net_19161_cascademuxed),
    .in3(net_19162),
    .lcout(net_15193),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_6 (
    .carryin(net_19158),
    .carryout(net_19164),
    .ce(),
    .clk(gnd),
    .in0(net_19165),
    .in1(net_19166),
    .in2(net_19167_cascademuxed),
    .in3(net_19168),
    .lcout(net_15194),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_2_7 (
    .carryin(net_19164),
    .carryout(net_19170),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19172),
    .in2(net_19173_cascademuxed),
    .in3(net_19174),
    .lcout(net_15195),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1000001000101000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_0 (
    .carryin(net_19214),
    .carryout(net_19251),
    .ce(),
    .clk(gnd),
    .in0(net_19252),
    .in1(net_19253),
    .in2(net_19254_cascademuxed),
    .in3(net_19255),
    .lcout(net_15347),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_1 (
    .carryin(net_19251),
    .carryout(net_19257),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19259),
    .in2(net_19260_cascademuxed),
    .in3(net_19261),
    .lcout(net_15348),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_2 (
    .carryin(net_19257),
    .carryout(net_19263),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19265),
    .in2(net_19266_cascademuxed),
    .in3(net_19267),
    .lcout(net_15349),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_3 (
    .carryin(net_19263),
    .carryout(net_19269),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19271),
    .in2(net_19272_cascademuxed),
    .in3(net_19273),
    .lcout(net_15350),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19276),
    .in1(net_19277),
    .in2(gnd),
    .in3(net_19279),
    .lcout(net_15351),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19298),
    .clk(net_19299),
    .in0(net_19282),
    .in1(net_19283),
    .in2(net_19284_cascademuxed),
    .in3(net_19285),
    .lcout(net_15352),
    .ltout(),
    .sr(net_19300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19298),
    .clk(net_19299),
    .in0(gnd),
    .in1(net_19289),
    .in2(net_19290_cascademuxed),
    .in3(net_19291),
    .lcout(net_15353),
    .ltout(),
    .sr(net_19300)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101001111110011),
    .SEQ_MODE(4'b0000)
  ) lc40_4_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19294),
    .in1(net_19295),
    .in2(net_19296_cascademuxed),
    .in3(net_19297),
    .lcout(net_15354),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111100001100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19422),
    .in0(gnd),
    .in1(net_19376),
    .in2(net_19377_cascademuxed),
    .in3(net_19378),
    .lcout(net_15470),
    .ltout(),
    .sr(net_19423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19422),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19384),
    .lcout(net_15471),
    .ltout(),
    .sr(net_19423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19422),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19390),
    .lcout(net_15472),
    .ltout(),
    .sr(net_19423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19422),
    .in0(net_19393),
    .in1(net_19394),
    .in2(net_19395_cascademuxed),
    .in3(net_19396),
    .lcout(net_15473),
    .ltout(),
    .sr(net_19423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000101010100000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19399),
    .in1(gnd),
    .in2(net_19401_cascademuxed),
    .in3(net_19402),
    .lcout(net_15474),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19422),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19408),
    .lcout(net_15475),
    .ltout(),
    .sr(net_19423)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19411),
    .in1(net_19412),
    .in2(net_19413_cascademuxed),
    .in3(net_19414),
    .lcout(net_15476),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(net_19498),
    .in1(gnd),
    .in2(net_19500_cascademuxed),
    .in3(gnd),
    .lcout(net_15593),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(gnd),
    .in1(net_19505),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15594),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19513),
    .lcout(net_15595),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_4_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19516),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19519),
    .lcout(net_15596),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19523),
    .in2(net_19524_cascademuxed),
    .in3(net_19525),
    .lcout(net_15597),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(gnd),
    .in1(net_19529),
    .in2(net_19530_cascademuxed),
    .in3(net_19531),
    .lcout(net_15598),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011101100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(net_19534),
    .in1(net_19535),
    .in2(net_19536_cascademuxed),
    .in3(net_19537),
    .lcout(net_15599),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_19545),
    .in0(gnd),
    .in1(net_19541),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15600),
    .ltout(),
    .sr(net_19546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19667),
    .clk(net_19668),
    .in0(gnd),
    .in1(gnd),
    .in2(net_19623_cascademuxed),
    .in3(gnd),
    .lcout(net_15716),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19627),
    .in1(gnd),
    .in2(net_19629_cascademuxed),
    .in3(gnd),
    .lcout(net_15717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19633),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19636),
    .lcout(net_15718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_19641_cascademuxed),
    .in3(net_19642),
    .lcout(net_15719),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101010001010),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19645),
    .in1(net_19646),
    .in2(net_19647_cascademuxed),
    .in3(net_19648),
    .lcout(net_15720),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19651),
    .in1(gnd),
    .in2(net_19653_cascademuxed),
    .in3(gnd),
    .lcout(net_15721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_19659_cascademuxed),
    .in3(net_19660),
    .lcout(net_15722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19667),
    .clk(net_19668),
    .in0(gnd),
    .in1(net_19664),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15723),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19744),
    .in1(net_19745),
    .in2(net_19746_cascademuxed),
    .in3(net_19747),
    .lcout(net_15839),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19790),
    .clk(net_19791),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_19753),
    .lcout(net_15840),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101001001010),
    .SEQ_MODE(4'b0000)
  ) lc40_4_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19756),
    .in1(net_19757),
    .in2(net_19758_cascademuxed),
    .in3(net_19759),
    .lcout(net_15841),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001000100010),
    .SEQ_MODE(4'b0000)
  ) lc40_4_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19762),
    .in1(net_19763),
    .in2(net_19764_cascademuxed),
    .in3(net_19765),
    .lcout(net_15842),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000001111),
    .SEQ_MODE(4'b0000)
  ) lc40_4_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_19768),
    .in1(net_19769),
    .in2(net_19770_cascademuxed),
    .in3(net_19771),
    .lcout(net_15843),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_4_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19790),
    .clk(net_19791),
    .in0(gnd),
    .in1(net_19775),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15844),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_4_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19790),
    .clk(net_19791),
    .in0(net_19780),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_15845),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_19790),
    .clk(net_19791),
    .in0(gnd),
    .in1(gnd),
    .in2(net_19788_cascademuxed),
    .in3(gnd),
    .lcout(net_15846),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_0 (
    .carryin(t175),
    .carryout(t177),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19868),
    .in2(net_19869_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_1 (
    .carryin(t177),
    .carryout(t178),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19874),
    .in2(net_19875_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_2 (
    .carryin(t178),
    .carryout(t179),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19880),
    .in2(net_19881_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_3 (
    .carryin(t179),
    .carryout(t180),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19886),
    .in2(net_19887_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_4 (
    .carryin(t180),
    .carryout(t181),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19892),
    .in2(net_19893_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_5 (
    .carryin(t181),
    .carryout(t182),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19898),
    .in2(net_19899_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_8_6 (
    .carryin(t182),
    .carryout(net_19902),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_19904),
    .in2(net_19905_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_8_7 (
    .carryin(net_19902),
    .carryout(net_19908),
    .ce(),
    .clk(net_19914),
    .in0(gnd),
    .in1(net_19910),
    .in2(net_19911_cascademuxed),
    .in3(net_19912),
    .lcout(net_15969),
    .ltout(),
    .sr(net_19915)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_0 (
    .carryin(net_19952),
    .carryout(net_19989),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_19991),
    .in2(net_19992_cascademuxed),
    .in3(net_19993),
    .lcout(net_16085),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_1 (
    .carryin(net_19989),
    .carryout(net_19995),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_19997),
    .in2(net_19998_cascademuxed),
    .in3(net_19999),
    .lcout(net_16086),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_2 (
    .carryin(net_19995),
    .carryout(net_20001),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20003),
    .in2(net_20004_cascademuxed),
    .in3(net_20005),
    .lcout(net_16087),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_3 (
    .carryin(net_20001),
    .carryout(net_20007),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20009),
    .in2(net_20010_cascademuxed),
    .in3(net_20011),
    .lcout(net_16088),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_4 (
    .carryin(net_20007),
    .carryout(net_20013),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20015),
    .in2(net_20016_cascademuxed),
    .in3(net_20017),
    .lcout(net_16089),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_5 (
    .carryin(net_20013),
    .carryout(net_20019),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20021),
    .in2(net_20022_cascademuxed),
    .in3(net_20023),
    .lcout(net_16090),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_6 (
    .carryin(net_20019),
    .carryout(net_20025),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20027),
    .in2(net_20028_cascademuxed),
    .in3(net_20029),
    .lcout(net_16091),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_9_7 (
    .carryin(net_20025),
    .carryout(net_20031),
    .ce(),
    .clk(net_20037),
    .in0(gnd),
    .in1(net_20033),
    .in2(net_20034_cascademuxed),
    .in3(net_20035),
    .lcout(net_16092),
    .ltout(),
    .sr(net_20038)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23947),
    .lcout(net_20039),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23953),
    .lcout(net_20040),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(net_23956),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20041),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23964_cascademuxed),
    .in3(gnd),
    .lcout(net_20042),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(net_23968),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20043),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(net_23974),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(gnd),
    .in1(net_23981),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23990),
    .clk(net_23991),
    .in0(net_23986),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(net_24067),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20162),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(net_24074),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20163),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24081_cascademuxed),
    .in3(gnd),
    .lcout(net_20164),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24087_cascademuxed),
    .in3(gnd),
    .lcout(net_20165),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(net_24092),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20166),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(net_24098),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20167),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(gnd),
    .in1(net_24104),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20168),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24114),
    .in0(net_24109),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20169),
    .ltout(),
    .sr(net_24115)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24193),
    .lcout(net_20285),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24199),
    .lcout(net_20286),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(net_24202),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20287),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24211),
    .lcout(net_20288),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24216_cascademuxed),
    .in3(gnd),
    .lcout(net_20289),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(net_24221),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20290),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(net_24226),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20291),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24237),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24235),
    .lcout(net_20292),
    .ltout(),
    .sr(net_24238)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(net_24313),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20408),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(net_24320),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20409),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24328),
    .lcout(net_20410),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24333_cascademuxed),
    .in3(gnd),
    .lcout(net_20411),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(net_24337),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20412),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(net_24344),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20413),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(net_24350),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20414),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24360),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24358),
    .lcout(net_20415),
    .ltout(),
    .sr(net_24361)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24438_cascademuxed),
    .in3(gnd),
    .lcout(net_20531),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(net_24443),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20532),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24451),
    .lcout(net_20533),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24462_cascademuxed),
    .in3(gnd),
    .lcout(net_20535),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24469),
    .lcout(net_20536),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24483),
    .in0(gnd),
    .in1(net_24479),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20538),
    .ltout(),
    .sr(net_24484)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(gnd),
    .in1(net_24566),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20655),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(net_24571),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20656),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(gnd),
    .in1(net_24578),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20657),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(net_24583),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20658),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(gnd),
    .in1(net_24590),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20659),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24598),
    .lcout(net_20660),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_24606),
    .in0(net_24601),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20661),
    .ltout(),
    .sr(net_24607)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24728),
    .clk(net_24729),
    .in0(net_24694),
    .in1(net_24695),
    .in2(net_24696_cascademuxed),
    .in3(net_24697),
    .lcout(net_20779),
    .ltout(),
    .sr(net_24730)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24728),
    .clk(net_24729),
    .in0(net_24712),
    .in1(net_24713),
    .in2(net_24714_cascademuxed),
    .in3(net_24715),
    .lcout(net_20782),
    .ltout(),
    .sr(net_24730)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24728),
    .clk(net_24729),
    .in0(net_24718),
    .in1(net_24719),
    .in2(net_24720_cascademuxed),
    .in3(net_24721),
    .lcout(net_20783),
    .ltout(),
    .sr(net_24730)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010111100000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24728),
    .clk(net_24729),
    .in0(net_24724),
    .in1(net_24725),
    .in2(net_24726_cascademuxed),
    .in3(net_24727),
    .lcout(net_20784),
    .ltout(),
    .sr(net_24730)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24851),
    .clk(net_24852),
    .in0(net_24811),
    .in1(net_24812),
    .in2(net_24813_cascademuxed),
    .in3(net_24814),
    .lcout(net_20901),
    .ltout(),
    .sr(net_24853)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24974),
    .clk(net_24975),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_24937),
    .lcout(net_21024),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_5_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_24948_cascademuxed),
    .in3(gnd),
    .lcout(net_21026),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_5_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_24952),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_21027),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_25098),
    .in0(gnd),
    .in1(gnd),
    .in2(net_25053_cascademuxed),
    .in3(gnd),
    .lcout(net_21146),
    .ltout(),
    .sr(net_25099)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_25098),
    .in0(gnd),
    .in1(gnd),
    .in2(net_25077_cascademuxed),
    .in3(gnd),
    .lcout(net_21150),
    .ltout(),
    .sr(net_25099)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_22844),
    .in0(net_22815),
    .in1(gnd),
    .in2(net_22817_cascademuxed),
    .in3(net_22818),
    .lcout(net_18894),
    .ltout(),
    .sr(net_22845)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_5_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_22841_cascademuxed),
    .in3(gnd),
    .lcout(net_18898),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23006),
    .clk(net_23007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_22968_cascademuxed),
    .in3(gnd),
    .lcout(net_19020),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23006),
    .clk(net_23007),
    .in0(net_22990),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19024),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_5_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_23095),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23129),
    .clk(net_23130),
    .in0(gnd),
    .in1(net_23108),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19182),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23129),
    .clk(net_23130),
    .in0(net_23113),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19183),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_5_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_23125),
    .in1(net_23126),
    .in2(net_23127_cascademuxed),
    .in3(net_23128),
    .lcout(net_19185),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(net_23206),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19301),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23215),
    .lcout(net_19302),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23220_cascademuxed),
    .in3(gnd),
    .lcout(net_19303),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(net_23224),
    .in1(net_23225),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19304),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23232_cascademuxed),
    .in3(gnd),
    .lcout(net_19305),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(net_23237),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19306),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(net_23243),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19307),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23253),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23251),
    .lcout(net_19308),
    .ltout(),
    .sr(net_23254)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_5_5_0 (
    .carryin(t264),
    .carryout(net_23328),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23330),
    .in2(net_23331_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_1 (
    .carryin(net_23328),
    .carryout(net_23334),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(net_23336),
    .in2(gnd),
    .in3(net_23338),
    .lcout(net_19425),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_2 (
    .carryin(net_23334),
    .carryout(net_23340),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(net_23342),
    .in2(gnd),
    .in3(net_23344),
    .lcout(net_19426),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_3 (
    .carryin(net_23340),
    .carryout(net_23346),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(net_23348),
    .in2(gnd),
    .in3(net_23350),
    .lcout(net_19427),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_4 (
    .carryin(net_23346),
    .carryout(net_23352),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(net_23354),
    .in2(gnd),
    .in3(net_23356),
    .lcout(net_19428),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_5 (
    .carryin(net_23352),
    .carryout(net_23358),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23361_cascademuxed),
    .in3(net_23362),
    .lcout(net_19429),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_6 (
    .carryin(net_23358),
    .carryout(net_23364),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(net_23366),
    .in2(gnd),
    .in3(net_23368),
    .lcout(net_19430),
    .ltout(),
    .sr(net_23377)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_5_5_7 (
    .carryin(net_23364),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23374),
    .lcout(net_19431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_0 (
    .carryin(t270),
    .carryout(net_23451),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23453),
    .in2(net_23454_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_1 (
    .carryin(net_23451),
    .carryout(net_23457),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23459),
    .in2(net_23460_cascademuxed),
    .in3(net_23461),
    .lcout(net_19548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_2 (
    .carryin(net_23457),
    .carryout(net_23463),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23465),
    .in2(net_23466_cascademuxed),
    .in3(net_23467),
    .lcout(net_19549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_3 (
    .carryin(net_23463),
    .carryout(net_23469),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23471),
    .in2(net_23472_cascademuxed),
    .in3(net_23473),
    .lcout(net_19550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_4 (
    .carryin(net_23469),
    .carryout(net_23475),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23477),
    .in2(net_23478_cascademuxed),
    .in3(net_23479),
    .lcout(net_19551),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_5 (
    .carryin(net_23475),
    .carryout(net_23481),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_23483),
    .in2(net_23484_cascademuxed),
    .in3(net_23485),
    .lcout(net_19552),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_5_6_6 (
    .carryin(net_23481),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23491),
    .lcout(net_19553),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23498),
    .clk(net_23499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23496_cascademuxed),
    .in3(gnd),
    .lcout(net_19554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101001001010),
    .SEQ_MODE(4'b0000)
  ) lc40_5_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_23581),
    .in1(net_23582),
    .in2(net_23583_cascademuxed),
    .in3(net_23584),
    .lcout(net_19671),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_23621),
    .clk(net_23622),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23589_cascademuxed),
    .in3(gnd),
    .lcout(net_19672),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000110010001100),
    .SEQ_MODE(4'b0000)
  ) lc40_5_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_23593),
    .in1(net_23594),
    .in2(net_23595_cascademuxed),
    .in3(gnd),
    .lcout(net_19673),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011011000100),
    .SEQ_MODE(4'b0000)
  ) lc40_5_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_23605),
    .in1(net_23606),
    .in2(net_23607_cascademuxed),
    .in3(net_23608),
    .lcout(net_19675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23700_cascademuxed),
    .in3(gnd),
    .lcout(net_19793),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(net_23704),
    .in1(gnd),
    .in2(net_23706_cascademuxed),
    .in3(gnd),
    .lcout(net_19794),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(gnd),
    .in1(net_23711),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19795),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110101010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(net_23716),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23719),
    .lcout(net_19796),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(net_23722),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19797),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(net_23728),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19798),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23736_cascademuxed),
    .in3(gnd),
    .lcout(net_19799),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23745),
    .in0(gnd),
    .in1(net_23741),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19800),
    .ltout(),
    .sr(net_23746)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(net_23822),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19916),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(net_23828),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19917),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(net_23834),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19918),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23842),
    .lcout(net_19919),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23848),
    .lcout(net_19920),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(net_23851),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_19921),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23860),
    .lcout(net_19922),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23868),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_23866),
    .lcout(net_19923),
    .ltout(),
    .sr(net_23869)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(net_30975),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27481),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30983_cascademuxed),
    .in3(gnd),
    .lcout(net_27482),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(gnd),
    .in1(net_30988),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27483),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(net_30993),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27484),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31001_cascademuxed),
    .in3(gnd),
    .lcout(net_27485),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(net_31011),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27487),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31022),
    .in0(gnd),
    .in1(net_31018),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27488),
    .ltout(),
    .sr(net_31023)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31100_cascademuxed),
    .in3(gnd),
    .lcout(net_27583),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(net_31104),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27584),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(gnd),
    .in1(net_31111),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27585),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(gnd),
    .in1(net_31117),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27586),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(gnd),
    .in1(net_31123),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27587),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(net_31128),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27588),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(net_31134),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27589),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31145),
    .in0(net_31140),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27590),
    .ltout(),
    .sr(net_31146)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_0 (
    .carryin(t383),
    .carryout(net_31220),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31222),
    .in2(net_31223_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_1 (
    .carryin(net_31220),
    .carryout(net_31226),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31228),
    .in2(net_31229_cascademuxed),
    .in3(net_31230),
    .lcout(net_27686),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_2 (
    .carryin(net_31226),
    .carryout(net_31232),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31234),
    .in2(net_31235_cascademuxed),
    .in3(net_31236),
    .lcout(net_27687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_3 (
    .carryin(net_31232),
    .carryout(net_31238),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31240),
    .in2(net_31241_cascademuxed),
    .in3(net_31242),
    .lcout(net_27688),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_4 (
    .carryin(net_31238),
    .carryout(net_31244),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31246),
    .in2(net_31247_cascademuxed),
    .in3(net_31248),
    .lcout(net_27689),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_5 (
    .carryin(net_31244),
    .carryout(net_31250),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31252),
    .in2(net_31253_cascademuxed),
    .in3(net_31254),
    .lcout(net_27690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_6 (
    .carryin(net_31250),
    .carryout(net_31256),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31258),
    .in2(net_31259_cascademuxed),
    .in3(net_31260),
    .lcout(net_27691),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_7 (
    .carryin(net_31256),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31266),
    .lcout(net_27692),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(net_31344),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27787),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31353),
    .lcout(net_27788),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(net_31356),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27789),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31364_cascademuxed),
    .in3(gnd),
    .lcout(net_27790),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(net_31368),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27791),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31376_cascademuxed),
    .in3(gnd),
    .lcout(net_27792),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31382_cascademuxed),
    .in3(gnd),
    .lcout(net_27793),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31391),
    .in0(net_31386),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27794),
    .ltout(),
    .sr(net_31392)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31514),
    .in0(gnd),
    .in1(net_31486),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27892),
    .ltout(),
    .sr(net_31515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31514),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31494),
    .lcout(net_27893),
    .ltout(),
    .sr(net_31515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31514),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31505_cascademuxed),
    .in3(gnd),
    .lcout(net_27895),
    .ltout(),
    .sr(net_31515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31514),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31511_cascademuxed),
    .in3(gnd),
    .lcout(net_27896),
    .ltout(),
    .sr(net_31515)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31590),
    .in1(net_31591),
    .in2(net_31592_cascademuxed),
    .in3(net_31593),
    .lcout(net_27991),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31596),
    .in1(net_31597),
    .in2(net_31598_cascademuxed),
    .in3(net_31599),
    .lcout(net_27992),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31602),
    .in1(net_31603),
    .in2(net_31604_cascademuxed),
    .in3(net_31605),
    .lcout(net_27993),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110010011000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31608),
    .in1(net_31609),
    .in2(net_31610_cascademuxed),
    .in3(net_31611),
    .lcout(net_27994),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31614),
    .in1(net_31615),
    .in2(net_31616_cascademuxed),
    .in3(net_31617),
    .lcout(net_27995),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010111100000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31620),
    .in1(net_31621),
    .in2(net_31622_cascademuxed),
    .in3(net_31623),
    .lcout(net_27996),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_7_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31628_cascademuxed),
    .in3(gnd),
    .lcout(net_27997),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010010100100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_31636),
    .clk(net_31637),
    .in0(net_31632),
    .in1(net_31633),
    .in2(net_31634_cascademuxed),
    .in3(net_31635),
    .lcout(net_27998),
    .ltout(),
    .sr(net_31638)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31760),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31716),
    .lcout(net_28093),
    .ltout(),
    .sr(net_31761)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31760),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31727_cascademuxed),
    .in3(gnd),
    .lcout(net_28095),
    .ltout(),
    .sr(net_31761)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31760),
    .in0(net_31731),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28096),
    .ltout(),
    .sr(net_31761)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31760),
    .in0(net_31737),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28097),
    .ltout(),
    .sr(net_31761)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31760),
    .in0(gnd),
    .in1(net_31756),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28100),
    .ltout(),
    .sr(net_31761)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_0 (
    .carryin(t442),
    .carryout(t445),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31837),
    .in2(net_31838_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_1 (
    .carryin(t445),
    .carryout(t447),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31843),
    .in2(net_31844_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_2 (
    .carryin(t447),
    .carryout(t449),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31849),
    .in2(net_31850_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_3 (
    .carryin(t449),
    .carryout(t451),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31855),
    .in2(net_31856_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_4 (
    .carryin(t451),
    .carryout(t453),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31861),
    .in2(net_31862_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_5 (
    .carryin(t453),
    .carryout(t455),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31867),
    .in2(net_31868_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_17_6 (
    .carryin(t455),
    .carryout(net_31871),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31873),
    .in2(net_31874_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011111111),
    .SEQ_MODE(4'b1000)
  ) lc40_7_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31883),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31881),
    .lcout(net_28202),
    .ltout(),
    .sr(net_31884)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_7_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31961_cascademuxed),
    .in3(gnd),
    .lcout(net_28297),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_7_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_31971),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28299),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_7_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31979_cascademuxed),
    .in3(gnd),
    .lcout(net_28300),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_32006),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31986),
    .lcout(net_28301),
    .ltout(),
    .sr(net_32007)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001111),
    .SEQ_MODE(4'b0000)
  ) lc40_7_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31991_cascademuxed),
    .in3(gnd),
    .lcout(net_28302),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_7_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_31995),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28303),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_32129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_32084_cascademuxed),
    .in3(gnd),
    .lcout(net_28399),
    .ltout(),
    .sr(net_32130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_32129),
    .in0(gnd),
    .in1(gnd),
    .in2(net_32102_cascademuxed),
    .in3(gnd),
    .lcout(net_28402),
    .ltout(),
    .sr(net_32130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_32129),
    .in0(gnd),
    .in1(net_32113),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28404),
    .ltout(),
    .sr(net_32130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_32129),
    .in0(gnd),
    .in1(net_32119),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_28405),
    .ltout(),
    .sr(net_32130)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_1_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_29875),
    .in0(net_29834),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26554),
    .ltout(),
    .sr(net_29876)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30038),
    .in0(net_30003),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26631),
    .ltout(),
    .sr(net_30039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30038),
    .in0(gnd),
    .in1(net_30010),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26632),
    .ltout(),
    .sr(net_30039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30038),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30018),
    .lcout(net_26633),
    .ltout(),
    .sr(net_30039)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30161),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30116_cascademuxed),
    .in3(gnd),
    .lcout(net_26767),
    .ltout(),
    .sr(net_30162)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30161),
    .in0(net_30126),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26769),
    .ltout(),
    .sr(net_30162)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30161),
    .in0(net_30132),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26770),
    .ltout(),
    .sr(net_30162)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30161),
    .in0(gnd),
    .in1(net_30139),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26771),
    .ltout(),
    .sr(net_30162)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(net_30237),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26869),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(gnd),
    .in1(net_30244),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26870),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30252),
    .lcout(net_26871),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(net_30255),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26872),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100000011000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(gnd),
    .in1(net_30268),
    .in2(net_30269_cascademuxed),
    .in3(gnd),
    .lcout(net_26874),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30284),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30281_cascademuxed),
    .in3(gnd),
    .lcout(net_26876),
    .ltout(),
    .sr(net_30285)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_0 (
    .carryin(t371),
    .carryout(net_30359),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_30361),
    .in2(net_30362_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_1 (
    .carryin(net_30359),
    .carryout(net_30365),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_30367),
    .in2(net_30368_cascademuxed),
    .in3(net_30369),
    .lcout(net_26972),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_2 (
    .carryin(net_30365),
    .carryout(net_30371),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_30373),
    .in2(net_30374_cascademuxed),
    .in3(net_30375),
    .lcout(net_26973),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_30378),
    .in1(gnd),
    .in2(net_30380_cascademuxed),
    .in3(net_30381),
    .lcout(net_26974),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111111100),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_30385),
    .in2(net_30386_cascademuxed),
    .in3(net_30387),
    .lcout(net_26975),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30392_cascademuxed),
    .in3(net_30393),
    .lcout(net_26976),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_30396),
    .in1(net_30397),
    .in2(net_30398_cascademuxed),
    .in3(net_30399),
    .lcout(net_26977),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30406),
    .clk(net_30407),
    .in0(gnd),
    .in1(net_30403),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_26978),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_6_0 (
    .carryin(t379),
    .carryout(net_30482),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_30484),
    .in2(net_30485_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_1 (
    .carryin(net_30482),
    .carryout(net_30488),
    .ce(),
    .clk(net_30530),
    .in0(gnd),
    .in1(net_30490),
    .in2(net_30491_cascademuxed),
    .in3(net_30492),
    .lcout(net_27074),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_2 (
    .carryin(net_30488),
    .carryout(net_30494),
    .ce(),
    .clk(net_30530),
    .in0(gnd),
    .in1(net_30496),
    .in2(net_30497_cascademuxed),
    .in3(net_30498),
    .lcout(net_27075),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30530),
    .in0(net_30501),
    .in1(net_30502),
    .in2(gnd),
    .in3(net_30504),
    .lcout(net_27076),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30530),
    .in0(gnd),
    .in1(net_30508),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27077),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30516),
    .lcout(net_27078),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30530),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30521_cascademuxed),
    .in3(gnd),
    .lcout(net_27079),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30530),
    .in0(net_30525),
    .in1(net_30526),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27080),
    .ltout(),
    .sr(net_30531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30608_cascademuxed),
    .in3(gnd),
    .lcout(net_27175),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30614_cascademuxed),
    .in3(gnd),
    .lcout(net_27176),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30621),
    .lcout(net_27177),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(net_30625),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27178),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(net_30630),
    .in1(gnd),
    .in2(net_30632_cascademuxed),
    .in3(gnd),
    .lcout(net_27179),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(net_30636),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30639),
    .lcout(net_27180),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30645),
    .lcout(net_27181),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30653),
    .in0(gnd),
    .in1(net_30649),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27182),
    .ltout(),
    .sr(net_30654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30732),
    .lcout(net_27277),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(net_30735),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27278),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30743_cascademuxed),
    .in3(gnd),
    .lcout(net_27279),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(net_30747),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27280),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30755_cascademuxed),
    .in3(gnd),
    .lcout(net_27281),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(net_30760),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27282),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(net_30766),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27283),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_30776),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30774),
    .lcout(net_27284),
    .ltout(),
    .sr(net_30777)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(net_30852),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27379),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30861),
    .lcout(net_27380),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(gnd),
    .in1(net_30865),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27381),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30873),
    .lcout(net_27382),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(net_30876),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_27383),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_30891),
    .lcout(net_27385),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_7_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_30898),
    .clk(net_30899),
    .in0(gnd),
    .in1(gnd),
    .in2(net_30896_cascademuxed),
    .in3(gnd),
    .lcout(net_27386),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34852),
    .clk(net_34853),
    .in0(gnd),
    .in1(net_34813),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30902),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34852),
    .clk(net_34853),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34820_cascademuxed),
    .in3(gnd),
    .lcout(net_30903),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34932),
    .lcout(net_31024),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34937_cascademuxed),
    .in3(gnd),
    .lcout(net_31025),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(gnd),
    .in1(net_34942),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31026),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(net_34947),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31027),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(net_34953),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31028),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34962),
    .lcout(net_31029),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34968),
    .lcout(net_31030),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34976),
    .in0(net_34971),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31031),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_0 (
    .carryin(t412),
    .carryout(t414),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_35053),
    .in2(net_35054_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_1 (
    .carryin(t414),
    .carryout(t415),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_35059),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_2 (
    .carryin(t415),
    .carryout(t416),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_35066_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_3 (
    .carryin(t416),
    .carryout(t417),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_35071),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_4 (
    .carryin(t417),
    .carryout(t418),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_35078_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_5 (
    .carryin(t418),
    .carryout(t419),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_35083),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_12_6 (
    .carryin(t419),
    .carryout(net_35087),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_35089),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_12_7 (
    .carryin(net_35087),
    .carryout(net_35093),
    .ce(),
    .clk(net_35099),
    .in0(gnd),
    .in1(net_35095),
    .in2(gnd),
    .in3(net_35097),
    .lcout(net_31154),
    .ltout(),
    .sr(net_35100)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_13_0 (
    .carryin(net_35137),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_35178),
    .lcout(net_31270),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(net_35181),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31271),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(gnd),
    .in1(gnd),
    .in2(net_35189_cascademuxed),
    .in3(gnd),
    .lcout(net_31272),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(net_35193),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31273),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_35202),
    .lcout(net_31274),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(gnd),
    .in1(gnd),
    .in2(net_35207_cascademuxed),
    .in3(gnd),
    .lcout(net_31275),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(gnd),
    .in1(net_35212),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31276),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35222),
    .in0(gnd),
    .in1(net_35218),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31277),
    .ltout(),
    .sr(net_35223)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35344),
    .clk(net_35345),
    .in0(net_35298),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_31393),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101111000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_35334),
    .in1(net_35335),
    .in2(net_35336_cascademuxed),
    .in3(net_35337),
    .lcout(net_31399),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35421),
    .in1(net_35422),
    .in2(net_35423_cascademuxed),
    .in3(net_35424),
    .lcout(net_31516),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35427),
    .in1(net_35428),
    .in2(net_35429_cascademuxed),
    .in3(net_35430),
    .lcout(net_31517),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35433),
    .in1(net_35434),
    .in2(net_35435_cascademuxed),
    .in3(net_35436),
    .lcout(net_31518),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010010100100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35439),
    .in1(net_35440),
    .in2(net_35441_cascademuxed),
    .in3(net_35442),
    .lcout(net_31519),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35445),
    .in1(net_35446),
    .in2(net_35447_cascademuxed),
    .in3(net_35448),
    .lcout(net_31520),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35457),
    .in1(net_35458),
    .in2(net_35459_cascademuxed),
    .in3(net_35460),
    .lcout(net_31522),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35467),
    .clk(net_35468),
    .in0(net_35463),
    .in1(net_35464),
    .in2(net_35465_cascademuxed),
    .in3(net_35466),
    .lcout(net_31523),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000011001010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35590),
    .clk(net_35591),
    .in0(net_35550),
    .in1(net_35551),
    .in2(net_35552_cascademuxed),
    .in3(net_35553),
    .lcout(net_31640),
    .ltout(),
    .sr(net_35592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35590),
    .clk(net_35591),
    .in0(net_35562),
    .in1(net_35563),
    .in2(net_35564_cascademuxed),
    .in3(net_35565),
    .lcout(net_31642),
    .ltout(),
    .sr(net_35592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101011011000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_35590),
    .clk(net_35591),
    .in0(net_35580),
    .in1(net_35581),
    .in2(net_35582_cascademuxed),
    .in3(net_35583),
    .lcout(net_31645),
    .ltout(),
    .sr(net_35592)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_1_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33706),
    .in0(gnd),
    .in1(gnd),
    .in2(net_33673_cascademuxed),
    .in3(gnd),
    .lcout(net_29755),
    .ltout(),
    .sr(net_33707)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33706),
    .in0(gnd),
    .in1(net_33678),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29756),
    .ltout(),
    .sr(net_33707)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_1_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33706),
    .in0(net_33689),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29758),
    .ltout(),
    .sr(net_33707)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33706),
    .in0(net_33695),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29759),
    .ltout(),
    .sr(net_33707)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33706),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_33704),
    .lcout(net_29760),
    .ltout(),
    .sr(net_33707)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33869),
    .in0(gnd),
    .in1(gnd),
    .in2(net_33824_cascademuxed),
    .in3(gnd),
    .lcout(net_29881),
    .ltout(),
    .sr(net_33870)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33869),
    .in0(gnd),
    .in1(net_33835),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29883),
    .ltout(),
    .sr(net_33870)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_33869),
    .in0(gnd),
    .in1(net_33859),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29887),
    .ltout(),
    .sr(net_33870)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110000101100),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33945),
    .in1(net_33946),
    .in2(net_33947_cascademuxed),
    .in3(net_33948),
    .lcout(net_30040),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_33991),
    .clk(net_33992),
    .in0(net_33975),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111110100000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33981),
    .in1(net_33982),
    .in2(net_33983_cascademuxed),
    .in3(net_33984),
    .lcout(net_30046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_33991),
    .clk(net_33992),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_33990),
    .lcout(net_30047),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34071),
    .lcout(net_30163),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(net_34080),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30165),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(net_34086),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30166),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(net_34092),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30167),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(gnd),
    .in1(net_34099),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30168),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34107),
    .lcout(net_30169),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34115),
    .in0(net_34110),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30170),
    .ltout(),
    .sr(net_34116)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(gnd),
    .in1(net_34192),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30286),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(net_34197),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30287),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34205_cascademuxed),
    .in3(gnd),
    .lcout(net_30288),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34212),
    .lcout(net_30289),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(net_34215),
    .in1(gnd),
    .in2(net_34217_cascademuxed),
    .in3(gnd),
    .lcout(net_30290),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(gnd),
    .in1(net_34222),
    .in2(gnd),
    .in3(net_34224),
    .lcout(net_30291),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(net_34227),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30292),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34238),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34235_cascademuxed),
    .in3(gnd),
    .lcout(net_30293),
    .ltout(),
    .sr(net_34239)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(net_34314),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30409),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34323),
    .lcout(net_30410),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(net_34332),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30412),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34341),
    .lcout(net_30413),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34346_cascademuxed),
    .in3(gnd),
    .lcout(net_30414),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34353),
    .lcout(net_30415),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_8_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34360),
    .clk(net_34361),
    .in0(net_34356),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30416),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34483),
    .clk(net_34484),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34439_cascademuxed),
    .in3(gnd),
    .lcout(net_30532),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34483),
    .clk(net_34484),
    .in0(gnd),
    .in1(net_34450),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30534),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34483),
    .clk(net_34484),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34476),
    .lcout(net_30538),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_0 (
    .carryin(t404),
    .carryout(net_34559),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34561),
    .in2(net_34562_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_1 (
    .carryin(net_34559),
    .carryout(net_34565),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34567),
    .in2(net_34568_cascademuxed),
    .in3(net_34569),
    .lcout(net_30656),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_2 (
    .carryin(net_34565),
    .carryout(net_34571),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34573),
    .in2(net_34574_cascademuxed),
    .in3(net_34575),
    .lcout(net_30657),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_3 (
    .carryin(net_34571),
    .carryout(net_34577),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34579),
    .in2(net_34580_cascademuxed),
    .in3(net_34581),
    .lcout(net_30658),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_4 (
    .carryin(net_34577),
    .carryout(net_34583),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34585),
    .in2(net_34586_cascademuxed),
    .in3(net_34587),
    .lcout(net_30659),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_5 (
    .carryin(net_34583),
    .carryout(net_34589),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34591),
    .in2(net_34592_cascademuxed),
    .in3(net_34593),
    .lcout(net_30660),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_6 (
    .carryin(net_34589),
    .carryout(net_34595),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34597),
    .in2(net_34598_cascademuxed),
    .in3(net_34599),
    .lcout(net_30661),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_8_7 (
    .carryin(net_34595),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34605),
    .lcout(net_30662),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34686),
    .lcout(net_30778),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_8_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34691_cascademuxed),
    .in3(net_34692),
    .lcout(net_30779),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(net_34696),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30780),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34709_cascademuxed),
    .in3(gnd),
    .lcout(net_30782),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(net_34714),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30783),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_34722),
    .lcout(net_30784),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34730),
    .in0(gnd),
    .in1(net_34726),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30785),
    .ltout(),
    .sr(net_34731)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38639_cascademuxed),
    .in3(gnd),
    .lcout(net_34732),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(net_38643),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34733),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(net_38649),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34734),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(gnd),
    .in1(net_38662),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34736),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38670),
    .lcout(net_34737),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38675_cascademuxed),
    .in3(gnd),
    .lcout(net_34738),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38684),
    .in0(net_38679),
    .in1(net_38680),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34739),
    .ltout(),
    .sr(net_38685)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000100010001),
    .SEQ_MODE(4'b1000)
  ) lc40_9_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38806),
    .clk(net_38807),
    .in0(net_38760),
    .in1(net_38761),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34855),
    .ltout(),
    .sr(net_38808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38806),
    .clk(net_38807),
    .in0(net_38796),
    .in1(net_38797),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34861),
    .ltout(),
    .sr(net_38808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38929),
    .clk(net_38930),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38886),
    .lcout(net_34978),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38929),
    .clk(net_38930),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38891_cascademuxed),
    .in3(gnd),
    .lcout(net_34979),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38929),
    .clk(net_38930),
    .in0(gnd),
    .in1(net_38908),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34982),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_38914),
    .in2(gnd),
    .in3(net_38916),
    .lcout(net_34983),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39052),
    .clk(net_39053),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39026_cascademuxed),
    .in3(gnd),
    .lcout(net_35104),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39052),
    .clk(net_39053),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_39039),
    .lcout(net_35106),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101100010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_9_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39042),
    .in1(net_39043),
    .in2(net_39044_cascademuxed),
    .in3(net_39045),
    .lcout(net_35107),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110011010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_9_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39129),
    .in1(net_39130),
    .in2(net_39131_cascademuxed),
    .in3(net_39132),
    .lcout(net_35224),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39175),
    .clk(net_39176),
    .in0(net_39141),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35226),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39175),
    .clk(net_39176),
    .in0(gnd),
    .in1(net_39148),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35227),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39175),
    .clk(net_39176),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_39156),
    .lcout(net_35228),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39175),
    .clk(net_39176),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_39162),
    .lcout(net_35229),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39175),
    .clk(net_39176),
    .in0(net_39171),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35231),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39254_cascademuxed),
    .in3(gnd),
    .lcout(net_35347),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110010001100),
    .SEQ_MODE(4'b0000)
  ) lc40_9_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39258),
    .in1(net_39259),
    .in2(net_39260_cascademuxed),
    .in3(net_39261),
    .lcout(net_35348),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39266_cascademuxed),
    .in3(gnd),
    .lcout(net_35349),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39272_cascademuxed),
    .in3(gnd),
    .lcout(net_35350),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39276),
    .in1(net_39277),
    .in2(net_39278_cascademuxed),
    .in3(net_39279),
    .lcout(net_35351),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39284_cascademuxed),
    .in3(gnd),
    .lcout(net_35352),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_39291),
    .lcout(net_35353),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39298),
    .clk(net_39299),
    .in0(net_39294),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35354),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39421),
    .clk(net_39422),
    .in0(gnd),
    .in1(net_39376),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35470),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39421),
    .clk(net_39422),
    .in0(gnd),
    .in1(net_39394),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35473),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39421),
    .clk(net_39422),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39401_cascademuxed),
    .in3(gnd),
    .lcout(net_35474),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39421),
    .clk(net_39422),
    .in0(gnd),
    .in1(net_39406),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35475),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39421),
    .clk(net_39422),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39419_cascademuxed),
    .in3(gnd),
    .lcout(net_35477),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39544),
    .clk(net_39545),
    .in0(net_39498),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_35593),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100001011000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39504),
    .in1(net_39505),
    .in2(net_39506_cascademuxed),
    .in3(net_39507),
    .lcout(net_35594),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_9_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_39510),
    .in1(net_39511),
    .in2(net_39512_cascademuxed),
    .in3(net_39513),
    .lcout(net_35595),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39544),
    .clk(net_39545),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39518_cascademuxed),
    .in3(gnd),
    .lcout(net_35596),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39621),
    .in1(net_39622),
    .in2(net_39623_cascademuxed),
    .in3(net_39624),
    .lcout(net_35716),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001011000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39627),
    .in1(net_39628),
    .in2(net_39629_cascademuxed),
    .in3(net_39630),
    .lcout(net_35717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39633),
    .in1(net_39634),
    .in2(net_39635_cascademuxed),
    .in3(net_39636),
    .lcout(net_35718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010010100100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39651),
    .in1(net_39652),
    .in2(net_39653_cascademuxed),
    .in3(net_39654),
    .lcout(net_35721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39657),
    .in1(net_39658),
    .in2(net_39659_cascademuxed),
    .in3(net_39660),
    .lcout(net_35722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101110010011000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(net_39663),
    .in1(net_39664),
    .in2(net_39665_cascademuxed),
    .in3(net_39666),
    .lcout(net_35723),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_1_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_37537),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37498_cascademuxed),
    .in3(gnd),
    .lcout(net_33585),
    .ltout(),
    .sr(net_37538)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_1_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_37537),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37510_cascademuxed),
    .in3(gnd),
    .lcout(net_33587),
    .ltout(),
    .sr(net_37538)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_1_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_37537),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37516_cascademuxed),
    .in3(gnd),
    .lcout(net_33588),
    .ltout(),
    .sr(net_37538)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_1_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_37537),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_37529),
    .lcout(net_33590),
    .ltout(),
    .sr(net_37538)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_37537),
    .in0(gnd),
    .in1(net_37533),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33591),
    .ltout(),
    .sr(net_37538)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37699),
    .clk(net_37700),
    .in0(gnd),
    .in1(net_37672),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33715),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37699),
    .clk(net_37700),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37691_cascademuxed),
    .in3(gnd),
    .lcout(net_33718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37822),
    .clk(net_37823),
    .in0(gnd),
    .in1(net_37795),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1101101010001010),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37812),
    .in1(net_37813),
    .in2(net_37814_cascademuxed),
    .in3(net_37815),
    .lcout(net_33877),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010110011110000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37899),
    .in1(net_37900),
    .in2(net_37901_cascademuxed),
    .in3(net_37902),
    .lcout(net_33994),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37945),
    .clk(net_37946),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_37914),
    .lcout(net_33996),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37945),
    .clk(net_37946),
    .in0(net_37929),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33999),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37945),
    .clk(net_37946),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37937_cascademuxed),
    .in3(gnd),
    .lcout(net_34000),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37945),
    .clk(net_37946),
    .in0(gnd),
    .in1(net_37942),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34001),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38024_cascademuxed),
    .in3(gnd),
    .lcout(net_34117),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38031),
    .lcout(net_34118),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(net_38040),
    .in1(net_38041),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34120),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(gnd),
    .in1(net_38047),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34121),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010000010100000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(net_38058),
    .in1(gnd),
    .in2(net_38060_cascademuxed),
    .in3(gnd),
    .lcout(net_34123),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38069),
    .in0(gnd),
    .in1(net_38065),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34124),
    .ltout(),
    .sr(net_38070)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38192),
    .in0(net_38145),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34240),
    .ltout(),
    .sr(net_38193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38192),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38160),
    .lcout(net_34242),
    .ltout(),
    .sr(net_38193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38192),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38166),
    .lcout(net_34243),
    .ltout(),
    .sr(net_38193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38192),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38172),
    .lcout(net_34244),
    .ltout(),
    .sr(net_38193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(gnd),
    .in1(net_38269),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34363),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38276_cascademuxed),
    .in3(gnd),
    .lcout(net_34364),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(net_38280),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34365),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(net_38286),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34366),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38294_cascademuxed),
    .in3(gnd),
    .lcout(net_34367),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000100010001000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(net_38298),
    .in1(net_38299),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34368),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(net_38304),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34369),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38315),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38312_cascademuxed),
    .in3(gnd),
    .lcout(net_34370),
    .ltout(),
    .sr(net_38316)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_0 (
    .carryin(t471),
    .carryout(net_38390),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_38392),
    .in2(net_38393_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_1 (
    .carryin(net_38390),
    .carryout(net_38396),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(net_38398),
    .in2(net_38399_cascademuxed),
    .in3(net_38400),
    .lcout(net_34487),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_2 (
    .carryin(net_38396),
    .carryout(net_38402),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(net_38404),
    .in2(gnd),
    .in3(net_38406),
    .lcout(net_34488),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_3 (
    .carryin(net_38402),
    .carryout(net_38408),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38411_cascademuxed),
    .in3(net_38412),
    .lcout(net_34489),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_4 (
    .carryin(net_38408),
    .carryout(net_38414),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(net_38416),
    .in2(gnd),
    .in3(net_38418),
    .lcout(net_34490),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_5 (
    .carryin(net_38414),
    .carryout(net_38420),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38423_cascademuxed),
    .in3(net_38424),
    .lcout(net_34491),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_6 (
    .carryin(net_38420),
    .carryout(net_38426),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38429_cascademuxed),
    .in3(net_38430),
    .lcout(net_34492),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_9_8_7 (
    .carryin(net_38426),
    .carryout(net_38432),
    .ce(),
    .clk(net_38438),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38435_cascademuxed),
    .in3(net_38436),
    .lcout(net_34493),
    .ltout(),
    .sr(net_38439)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b1111111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_9_0 (
    .carryin(net_38476),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38517),
    .lcout(net_34609),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38522_cascademuxed),
    .in3(gnd),
    .lcout(net_34610),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38528_cascademuxed),
    .in3(gnd),
    .lcout(net_34611),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(net_38532),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34612),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(gnd),
    .in1(net_38539),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34613),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(net_38544),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34614),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(net_38550),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34615),
    .ltout(),
    .sr(net_38562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_38561),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38559),
    .lcout(net_34616),
    .ltout(),
    .sr(net_38562)
  );
  Odrv4 odrv_0_10_2158_1656 (
    .I(net_2158),
    .O(net_1656)
  );
  Odrv4 odrv_0_10_2159_1658 (
    .I(net_2159),
    .O(net_1658)
  );
  Odrv4 odrv_0_10_2160_2287 (
    .I(net_2160),
    .O(net_2287)
  );
  Odrv4 odrv_0_10_2161_2289 (
    .I(net_2161),
    .O(net_2289)
  );
  Odrv4 odrv_0_10_2162_2273 (
    .I(net_2162),
    .O(net_2273)
  );
  Odrv4 odrv_0_10_2163_2293 (
    .I(net_2163),
    .O(net_2293)
  );
  Odrv4 odrv_0_10_2164_2295 (
    .I(net_2164),
    .O(net_2295)
  );
  Odrv4 odrv_0_10_2165_2297 (
    .I(net_2165),
    .O(net_2297)
  );
  Odrv4 odrv_0_11_2364_2478 (
    .I(net_2364),
    .O(net_2478)
  );
  Odrv4 odrv_0_11_2365_2488 (
    .I(net_2365),
    .O(net_2488)
  );
  Odrv4 odrv_0_11_2366_2490 (
    .I(net_2366),
    .O(net_2490)
  );
  Odrv4 odrv_0_11_2367_2446 (
    .I(net_2367),
    .O(net_2446)
  );
  Odrv4 odrv_0_11_2368_2448 (
    .I(net_2368),
    .O(net_2448)
  );
  Odrv4 odrv_0_11_2369_2485 (
    .I(net_2369),
    .O(net_2485)
  );
  Odrv4 odrv_0_11_2370_2444 (
    .I(net_2370),
    .O(net_2444)
  );
  Odrv4 odrv_0_11_2371_2456 (
    .I(net_2371),
    .O(net_2456)
  );
  Odrv4 odrv_0_12_2572_2660 (
    .I(net_2572),
    .O(net_2660)
  );
  Odrv4 odrv_0_12_2573_2309 (
    .I(net_2573),
    .O(net_2309)
  );
  Odrv4 odrv_0_12_2574_2665 (
    .I(net_2574),
    .O(net_2665)
  );
  Odrv4 odrv_0_12_2575_2703 (
    .I(net_2575),
    .O(net_2703)
  );
  Odrv4 odrv_0_12_2576_2492 (
    .I(net_2576),
    .O(net_2492)
  );
  Odrv4 odrv_0_12_2577_2086 (
    .I(net_2577),
    .O(net_2086)
  );
  Odrv4 odrv_0_12_2578_2088 (
    .I(net_2578),
    .O(net_2088)
  );
  Odrv4 odrv_0_12_2579_2498 (
    .I(net_2579),
    .O(net_2498)
  );
  Odrv4 odrv_0_13_2781_2861 (
    .I(net_2781),
    .O(net_2861)
  );
  Odrv4 odrv_0_13_2782_2288 (
    .I(net_2782),
    .O(net_2288)
  );
  Odrv4 odrv_0_13_2783_2501 (
    .I(net_2783),
    .O(net_2501)
  );
  Odrv4 odrv_0_13_2784_2893 (
    .I(net_2784),
    .O(net_2893)
  );
  Odrv4 odrv_0_13_2785_2878 (
    .I(net_2785),
    .O(net_2878)
  );
  Odrv4 odrv_0_13_2786_2702 (
    .I(net_2786),
    .O(net_2702)
  );
  Odrv4 odrv_0_13_2787_2298 (
    .I(net_2787),
    .O(net_2298)
  );
  Odrv4 odrv_0_15_3218_3306 (
    .I(net_3218),
    .O(net_3306)
  );
  Odrv4 odrv_0_15_3219_3308 (
    .I(net_3219),
    .O(net_3308)
  );
  Odrv4 odrv_0_15_3220_2720 (
    .I(net_3220),
    .O(net_2720)
  );
  Odrv4 odrv_0_15_3221_2920 (
    .I(net_3221),
    .O(net_2920)
  );
  Odrv4 odrv_0_15_3222_3344 (
    .I(net_3222),
    .O(net_3344)
  );
  Odrv4 odrv_0_15_3223_3300 (
    .I(net_3223),
    .O(net_3300)
  );
  Odrv4 odrv_0_15_3224_2926 (
    .I(net_3224),
    .O(net_2926)
  );
  Odrv4 odrv_0_15_3225_3304 (
    .I(net_3225),
    .O(net_3304)
  );
  Odrv4 odrv_0_16_3424_2913 (
    .I(net_3424),
    .O(net_2913)
  );
  Odrv4 odrv_0_16_3425_2719 (
    .I(net_3425),
    .O(net_2719)
  );
  Odrv4 odrv_0_16_3426_2721 (
    .I(net_3426),
    .O(net_2721)
  );
  Odrv4 odrv_0_16_3427_3151 (
    .I(net_3427),
    .O(net_3151)
  );
  Odrv4 odrv_0_16_3428_3137 (
    .I(net_3428),
    .O(net_3137)
  );
  Odrv4 odrv_0_16_3429_3139 (
    .I(net_3429),
    .O(net_3139)
  );
  Odrv4 odrv_0_16_3430_3157 (
    .I(net_3430),
    .O(net_3157)
  );
  Odrv4 odrv_0_16_3431_3514 (
    .I(net_3431),
    .O(net_3514)
  );
  Odrv4 odrv_0_17_3632_3351 (
    .I(net_3632),
    .O(net_3351)
  );
  Odrv4 odrv_0_17_3633_3562 (
    .I(net_3633),
    .O(net_3562)
  );
  Odrv4 odrv_0_17_3634_3746 (
    .I(net_3634),
    .O(net_3746)
  );
  Odrv4 odrv_0_17_3635_3158 (
    .I(net_3635),
    .O(net_3158)
  );
  Odrv4 odrv_0_17_3636_3758 (
    .I(net_3636),
    .O(net_3758)
  );
  Odrv4 odrv_0_17_3637_3731 (
    .I(net_3637),
    .O(net_3731)
  );
  Odrv4 odrv_0_17_3638_3556 (
    .I(net_3638),
    .O(net_3556)
  );
  Odrv4 odrv_0_17_3639_3365 (
    .I(net_3639),
    .O(net_3365)
  );
  Odrv4 odrv_0_18_3841_3362 (
    .I(net_3841),
    .O(net_3362)
  );
  Odrv4 odrv_0_18_3842_3559 (
    .I(net_3842),
    .O(net_3559)
  );
  Odrv4 odrv_0_18_3843_3350 (
    .I(net_3843),
    .O(net_3350)
  );
  Odrv4 odrv_0_18_3844_3965 (
    .I(net_3844),
    .O(net_3965)
  );
  Odrv4 odrv_0_18_3845_3354 (
    .I(net_3845),
    .O(net_3354)
  );
  Odrv4 odrv_0_18_3846_3356 (
    .I(net_3846),
    .O(net_3356)
  );
  Odrv4 odrv_0_18_3847_3553 (
    .I(net_3847),
    .O(net_3553)
  );
  Odrv4 odrv_0_23_4959_5039 (
    .I(net_4959),
    .O(net_5039)
  );
  Odrv4 odrv_0_23_4960_4425 (
    .I(net_4960),
    .O(net_4425)
  );
  Odrv4 odrv_0_23_4961_4427 (
    .I(net_4961),
    .O(net_4427)
  );
  Odrv4 odrv_0_23_4962_4429 (
    .I(net_4962),
    .O(net_4429)
  );
  Odrv4 odrv_0_23_4963_4431 (
    .I(net_4963),
    .O(net_4431)
  );
  Odrv4 odrv_0_23_4964_4433 (
    .I(net_4964),
    .O(net_4433)
  );
  Odrv4 odrv_0_23_4965_4435 (
    .I(net_4965),
    .O(net_4435)
  );
  Odrv4 odrv_0_23_4966_4653 (
    .I(net_4966),
    .O(net_4653)
  );
  Odrv4 odrv_0_24_5165_4654 (
    .I(net_5165),
    .O(net_4654)
  );
  Odrv4 odrv_0_24_5166_5260 (
    .I(net_5166),
    .O(net_5260)
  );
  Odrv4 odrv_0_24_5167_4658 (
    .I(net_5167),
    .O(net_4658)
  );
  Odrv4 odrv_0_24_5168_4660 (
    .I(net_5168),
    .O(net_4660)
  );
  Odrv4 odrv_0_24_5169_5091 (
    .I(net_5169),
    .O(net_5091)
  );
  Odrv4 odrv_0_24_5170_4880 (
    .I(net_5170),
    .O(net_4880)
  );
  Odrv4 odrv_0_24_5171_4650 (
    .I(net_5171),
    .O(net_4650)
  );
  Odrv4 odrv_0_24_5172_5097 (
    .I(net_5172),
    .O(net_5097)
  );
  Odrv4 odrv_0_25_5373_5453 (
    .I(net_5373),
    .O(net_5453)
  );
  Odrv4 odrv_0_25_5374_4879 (
    .I(net_5374),
    .O(net_4879)
  );
  Odrv4 odrv_0_25_5375_4881 (
    .I(net_5375),
    .O(net_4881)
  );
  Odrv4 odrv_0_25_5376_5497 (
    .I(net_5376),
    .O(net_5497)
  );
  Odrv4 odrv_0_25_5377_5499 (
    .I(net_5377),
    .O(net_5499)
  );
  Odrv4 odrv_0_25_5378_5472 (
    .I(net_5378),
    .O(net_5472)
  );
  Odrv4 odrv_0_25_5379_5088 (
    .I(net_5379),
    .O(net_5088)
  );
  Odrv4 odrv_0_25_5380_5299 (
    .I(net_5380),
    .O(net_5299)
  );
  Odrv4 odrv_0_26_5582_5298 (
    .I(net_5582),
    .O(net_5298)
  );
  Odrv4 odrv_0_26_5583_5511 (
    .I(net_5583),
    .O(net_5511)
  );
  Odrv4 odrv_0_26_5584_5302 (
    .I(net_5584),
    .O(net_5302)
  );
  Odrv4 odrv_0_26_5585_5093 (
    .I(net_5585),
    .O(net_5093)
  );
  Odrv4 odrv_0_26_5586_5095 (
    .I(net_5586),
    .O(net_5095)
  );
  Odrv4 odrv_0_26_5587_4900 (
    .I(net_5587),
    .O(net_4900)
  );
  Odrv4 odrv_0_26_5588_5683 (
    .I(net_5588),
    .O(net_5683)
  );
  Odrv4 odrv_0_5_1098_1178 (
    .I(net_1098),
    .O(net_1178)
  );
  Odrv4 odrv_0_5_1099_1206 (
    .I(net_1099),
    .O(net_1206)
  );
  Odrv4 odrv_0_5_1100_798 (
    .I(net_1100),
    .O(net_798)
  );
  Odrv4 odrv_0_5_1101_1210 (
    .I(net_1101),
    .O(net_1210)
  );
  Odrv4 odrv_0_5_1102_1195 (
    .I(net_1102),
    .O(net_1195)
  );
  Odrv4 odrv_0_5_1103_804 (
    .I(net_1103),
    .O(net_804)
  );
  Odrv4 odrv_0_5_1104_1199 (
    .I(net_1104),
    .O(net_1199)
  );
  Odrv4 odrv_0_5_1105_1184 (
    .I(net_1105),
    .O(net_1184)
  );
  Odrv4 odrv_0_6_1304_1418 (
    .I(net_1304),
    .O(net_1418)
  );
  Odrv4 odrv_0_6_1305_811 (
    .I(net_1305),
    .O(net_811)
  );
  Odrv4 odrv_0_6_1306_1430 (
    .I(net_1306),
    .O(net_1430)
  );
  Odrv4 odrv_0_6_1307_1228 (
    .I(net_1307),
    .O(net_1228)
  );
  Odrv4 odrv_0_6_1308_1423 (
    .I(net_1308),
    .O(net_1423)
  );
  Odrv4 odrv_0_6_1309_1019 (
    .I(net_1309),
    .O(net_1019)
  );
  Odrv4 odrv_0_6_1310_1384 (
    .I(net_1310),
    .O(net_1384)
  );
  Odrv4 odrv_0_6_1311_1023 (
    .I(net_1311),
    .O(net_1023)
  );
  Odrv4 odrv_0_7_1512_1618 (
    .I(net_1512),
    .O(net_1618)
  );
  Odrv4 odrv_0_7_1513_1233 (
    .I(net_1513),
    .O(net_1233)
  );
  Odrv4 odrv_0_7_1514_1235 (
    .I(net_1514),
    .O(net_1235)
  );
  Odrv4 odrv_0_7_1515_1636 (
    .I(net_1515),
    .O(net_1636)
  );
  Odrv4 odrv_0_7_1516_1645 (
    .I(net_1516),
    .O(net_1645)
  );
  Odrv4 odrv_0_7_1517_1594 (
    .I(net_1517),
    .O(net_1594)
  );
  Odrv4 odrv_0_7_1518_1227 (
    .I(net_1518),
    .O(net_1227)
  );
  Odrv4 odrv_0_7_1519_1598 (
    .I(net_1519),
    .O(net_1598)
  );
  Odrv4 odrv_0_8_1721_1801 (
    .I(net_1721),
    .O(net_1801)
  );
  Odrv4 odrv_0_8_1722_1031 (
    .I(net_1722),
    .O(net_1031)
  );
  Odrv4 odrv_0_8_1723_1814 (
    .I(net_1723),
    .O(net_1814)
  );
  Odrv4 odrv_0_8_1724_1232 (
    .I(net_1724),
    .O(net_1232)
  );
  Odrv4 odrv_0_8_1725_1037 (
    .I(net_1725),
    .O(net_1037)
  );
  Odrv4 odrv_0_8_1726_1447 (
    .I(net_1726),
    .O(net_1447)
  );
  Odrv4 odrv_0_8_1727_1805 (
    .I(net_1727),
    .O(net_1805)
  );
  Odrv4 odrv_10_10_38563_34877 (
    .I(net_38563),
    .O(net_34877)
  );
  Odrv4 odrv_10_10_38563_38596 (
    .I(net_38563),
    .O(net_38596)
  );
  Odrv4 odrv_10_10_38563_42529 (
    .I(net_38563),
    .O(net_42529)
  );
  Odrv4 odrv_10_10_38565_38346 (
    .I(net_38565),
    .O(net_38346)
  );
  Odrv12 odrv_10_10_38569_2200 (
    .I(net_38569),
    .O(net_2200)
  );
  Odrv4 odrv_10_10_38569_34873 (
    .I(net_38569),
    .O(net_34873)
  );
  Odrv4 odrv_10_10_38570_38466 (
    .I(net_38570),
    .O(net_38466)
  );
  Odrv4 odrv_10_10_38570_38703 (
    .I(net_38570),
    .O(net_38703)
  );
  Odrv4 odrv_10_10_38570_38720 (
    .I(net_38570),
    .O(net_38720)
  );
  Odrv4 odrv_10_11_38690_34990 (
    .I(net_38690),
    .O(net_34990)
  );
  Odrv4 odrv_10_11_38693_34998 (
    .I(net_38693),
    .O(net_34998)
  );
  Odrv4 odrv_10_12_38811_38955 (
    .I(net_38811),
    .O(net_38955)
  );
  Odrv4 odrv_10_14_39055_39197 (
    .I(net_39055),
    .O(net_39197)
  );
  Odrv4 odrv_10_14_39056_42794 (
    .I(net_39056),
    .O(net_42794)
  );
  Odrv4 odrv_10_14_39058_42798 (
    .I(net_39058),
    .O(net_42798)
  );
  Odrv4 odrv_10_14_39059_35359 (
    .I(net_39059),
    .O(net_35359)
  );
  Odrv4 odrv_10_14_39060_43023 (
    .I(net_39060),
    .O(net_43023)
  );
  Odrv4 odrv_10_14_39062_38958 (
    .I(net_39062),
    .O(net_38958)
  );
  Odrv4 odrv_10_15_39180_39325 (
    .I(net_39180),
    .O(net_39325)
  );
  Odrv4 odrv_10_18_39547_43513 (
    .I(net_39547),
    .O(net_43513)
  );
  Odrv4 odrv_10_18_39551_43523 (
    .I(net_39551),
    .O(net_43523)
  );
  Odrv4 odrv_10_19_39671_43281 (
    .I(net_39671),
    .O(net_43281)
  );
  Odrv4 odrv_10_19_39677_43405 (
    .I(net_39677),
    .O(net_43405)
  );
  Odrv4 odrv_10_1_37422_41440 (
    .I(net_37422),
    .O(net_41440)
  );
  Odrv4 odrv_10_3_37708_37597 (
    .I(net_37708),
    .O(net_37597)
  );
  Odrv12 odrv_10_4_37825_41270 (
    .I(net_37825),
    .O(net_41270)
  );
  Odrv4 odrv_10_4_37830_41793 (
    .I(net_37830),
    .O(net_41793)
  );
  Odrv4 odrv_10_4_37832_41686 (
    .I(net_37832),
    .O(net_41686)
  );
  Odrv4 odrv_10_5_37949_37729 (
    .I(net_37949),
    .O(net_37729)
  );
  Odrv4 odrv_10_5_37954_37849 (
    .I(net_37954),
    .O(net_37849)
  );
  Odrv4 odrv_10_6_38072_42041 (
    .I(net_38072),
    .O(net_42041)
  );
  Odrv4 odrv_10_6_38075_34375 (
    .I(net_38075),
    .O(net_34375)
  );
  Odrv4 odrv_10_6_38078_38102 (
    .I(net_38078),
    .O(net_38102)
  );
  Odrv4 odrv_10_7_38194_38336 (
    .I(net_38194),
    .O(net_38336)
  );
  Odrv4 odrv_10_7_38194_42057 (
    .I(net_38194),
    .O(net_42057)
  );
  Odrv4 odrv_10_7_38198_34498 (
    .I(net_38198),
    .O(net_34498)
  );
  Odrv4 odrv_10_7_38198_38219 (
    .I(net_38198),
    .O(net_38219)
  );
  Odrv4 odrv_10_7_38199_37983 (
    .I(net_38199),
    .O(net_37983)
  );
  Odrv4 odrv_10_8_38317_41926 (
    .I(net_38317),
    .O(net_41926)
  );
  Odrv4 odrv_10_8_38324_30793 (
    .I(net_38324),
    .O(net_30793)
  );
  Odrv4 odrv_10_8_38324_38457 (
    .I(net_38324),
    .O(net_38457)
  );
  Odrv4 odrv_10_8_38324_42306 (
    .I(net_38324),
    .O(net_42306)
  );
  Odrv12 odrv_10_9_38443_42281 (
    .I(net_38443),
    .O(net_42281)
  );
  Odrv4 odrv_11_11_42517_42659 (
    .I(net_42517),
    .O(net_42659)
  );
  Odrv12 odrv_11_11_42519_45216 (
    .I(net_42519),
    .O(net_45216)
  );
  Odrv4 odrv_11_11_42519_46258 (
    .I(net_42519),
    .O(net_46258)
  );
  Odrv4 odrv_11_11_42520_46260 (
    .I(net_42520),
    .O(net_46260)
  );
  Odrv12 odrv_11_11_42520_46358 (
    .I(net_42520),
    .O(net_46358)
  );
  Odrv12 odrv_11_11_42524_2407 (
    .I(net_42524),
    .O(net_2407)
  );
  Odrv4 odrv_11_11_42524_46252 (
    .I(net_42524),
    .O(net_46252)
  );
  Odrv4 odrv_11_12_42640_46249 (
    .I(net_42640),
    .O(net_46249)
  );
  Odrv4 odrv_11_12_42641_46610 (
    .I(net_42641),
    .O(net_46610)
  );
  Odrv4 odrv_11_12_42644_42791 (
    .I(net_42644),
    .O(net_42791)
  );
  Odrv12 odrv_11_12_42645_45743 (
    .I(net_42645),
    .O(net_45743)
  );
  Odrv4 odrv_11_13_42765_42672 (
    .I(net_42765),
    .O(net_42672)
  );
  Odrv4 odrv_11_14_42886_46852 (
    .I(net_42886),
    .O(net_46852)
  );
  Odrv4 odrv_11_14_42888_46627 (
    .I(net_42888),
    .O(net_46627)
  );
  Odrv12 odrv_11_14_42890_45867 (
    .I(net_42890),
    .O(net_45867)
  );
  Odrv4 odrv_11_14_42891_35368 (
    .I(net_42891),
    .O(net_35368)
  );
  Odrv12 odrv_11_14_42893_46235 (
    .I(net_42893),
    .O(net_46235)
  );
  Odrv4 odrv_11_15_43010_43044 (
    .I(net_43010),
    .O(net_43044)
  );
  Odrv4 odrv_11_15_43011_43156 (
    .I(net_43011),
    .O(net_43156)
  );
  Odrv4 odrv_11_15_43013_43034 (
    .I(net_43013),
    .O(net_43034)
  );
  Odrv4 odrv_11_15_43016_35485 (
    .I(net_43016),
    .O(net_35485)
  );
  Odrv4 odrv_11_16_43132_43165 (
    .I(net_43132),
    .O(net_43165)
  );
  Odrv4 odrv_11_16_43133_43276 (
    .I(net_43133),
    .O(net_43276)
  );
  Odrv4 odrv_11_18_43380_47119 (
    .I(net_43380),
    .O(net_47119)
  );
  Odrv4 odrv_11_18_43383_47235 (
    .I(net_43383),
    .O(net_47235)
  );
  Odrv4 odrv_11_18_43385_47113 (
    .I(net_43385),
    .O(net_47113)
  );
  Odrv4 odrv_11_1_41250_45276 (
    .I(net_41250),
    .O(net_45276)
  );
  Odrv4 odrv_11_2_41375_37716 (
    .I(net_41375),
    .O(net_37716)
  );
  Odrv4 odrv_11_2_41379_45378 (
    .I(net_41379),
    .O(net_45378)
  );
  Odrv4 odrv_11_2_41380_37720 (
    .I(net_41380),
    .O(net_37720)
  );
  Odrv4 odrv_11_4_41657_41431 (
    .I(net_41657),
    .O(net_41431)
  );
  Odrv4 odrv_11_4_41658_45264 (
    .I(net_41658),
    .O(net_45264)
  );
  Odrv4 odrv_11_4_41660_45632 (
    .I(net_41660),
    .O(net_45632)
  );
  Odrv4 odrv_11_4_41662_37966 (
    .I(net_41662),
    .O(net_37966)
  );
  Odrv12 odrv_11_4_41663_34126 (
    .I(net_41663),
    .O(net_34126)
  );
  Odrv4 odrv_11_4_41663_41559 (
    .I(net_41663),
    .O(net_41559)
  );
  Odrv4 odrv_11_5_41779_41558 (
    .I(net_41779),
    .O(net_41558)
  );
  Odrv4 odrv_11_5_41780_41560 (
    .I(net_41780),
    .O(net_41560)
  );
  Odrv4 odrv_11_5_41781_41688 (
    .I(net_41781),
    .O(net_41688)
  );
  Odrv4 odrv_11_5_41781_45751 (
    .I(net_41781),
    .O(net_45751)
  );
  Odrv4 odrv_11_5_41782_41564 (
    .I(net_41782),
    .O(net_41564)
  );
  Odrv4 odrv_11_5_41783_41566 (
    .I(net_41783),
    .O(net_41566)
  );
  Odrv4 odrv_11_5_41784_38087 (
    .I(net_41784),
    .O(net_38087)
  );
  Odrv4 odrv_11_5_41784_45747 (
    .I(net_41784),
    .O(net_45747)
  );
  Odrv4 odrv_11_5_41784_45764 (
    .I(net_41784),
    .O(net_45764)
  );
  Odrv4 odrv_11_5_41786_41682 (
    .I(net_41786),
    .O(net_41682)
  );
  Odrv4 odrv_11_6_41903_42046 (
    .I(net_41903),
    .O(net_42046)
  );
  Odrv4 odrv_11_6_41903_45767 (
    .I(net_41903),
    .O(net_45767)
  );
  Odrv4 odrv_11_6_41903_45872 (
    .I(net_41903),
    .O(net_45872)
  );
  Odrv4 odrv_11_7_42025_45991 (
    .I(net_42025),
    .O(net_45991)
  );
  Odrv4 odrv_11_7_42029_46008 (
    .I(net_42029),
    .O(net_46008)
  );
  Odrv4 odrv_11_7_42030_45993 (
    .I(net_42030),
    .O(net_45993)
  );
  Odrv4 odrv_11_8_42148_45885 (
    .I(net_42148),
    .O(net_45885)
  );
  Odrv4 odrv_11_8_42148_46011 (
    .I(net_42148),
    .O(net_46011)
  );
  Odrv4 odrv_11_8_42150_41931 (
    .I(net_42150),
    .O(net_41931)
  );
  Odrv4 odrv_11_8_42150_42294 (
    .I(net_42150),
    .O(net_42294)
  );
  Odrv4 odrv_11_8_42150_45889 (
    .I(net_42150),
    .O(net_45889)
  );
  Odrv12 odrv_11_8_42151_19925 (
    .I(net_42151),
    .O(net_19925)
  );
  Odrv4 odrv_11_8_42151_34626 (
    .I(net_42151),
    .O(net_34626)
  );
  Odrv4 odrv_11_8_42153_34630 (
    .I(net_42153),
    .O(net_34630)
  );
  Odrv12 odrv_11_8_42153_45215 (
    .I(net_42153),
    .O(net_45215)
  );
  Odrv4 odrv_11_8_42154_34632 (
    .I(net_42154),
    .O(net_34632)
  );
  Odrv12 odrv_11_8_42154_7898 (
    .I(net_42154),
    .O(net_7898)
  );
  Odrv12 odrv_11_8_42155_1764 (
    .I(net_42155),
    .O(net_1764)
  );
  Odrv4 odrv_11_8_42155_34624 (
    .I(net_42155),
    .O(net_34624)
  );
  Odrv4 odrv_11_9_42275_42296 (
    .I(net_42275),
    .O(net_42296)
  );
  Odrv4 odrv_11_9_42278_42302 (
    .I(net_42278),
    .O(net_42302)
  );
  Odrv4 odrv_12_10_46226_46132 (
    .I(net_46226),
    .O(net_46132)
  );
  Odrv4 odrv_12_10_46226_46369 (
    .I(net_46226),
    .O(net_46369)
  );
  Odrv4 odrv_12_10_46228_50206 (
    .I(net_46228),
    .O(net_50206)
  );
  Odrv4 odrv_12_10_46229_46012 (
    .I(net_46229),
    .O(net_46012)
  );
  Odrv4 odrv_12_10_46229_46250 (
    .I(net_46229),
    .O(net_46250)
  );
  Odrv4 odrv_12_10_46229_46376 (
    .I(net_46229),
    .O(net_46376)
  );
  Odrv4 odrv_12_10_46231_50212 (
    .I(net_46231),
    .O(net_50212)
  );
  Odrv4 odrv_12_10_46232_38701 (
    .I(net_46232),
    .O(net_38701)
  );
  Odrv4 odrv_12_10_46232_46365 (
    .I(net_46232),
    .O(net_46365)
  );
  Odrv4 odrv_12_10_46232_50086 (
    .I(net_46232),
    .O(net_50086)
  );
  Odrv4 odrv_12_10_46232_50214 (
    .I(net_46232),
    .O(net_50214)
  );
  Odrv4 odrv_12_11_46350_50320 (
    .I(net_46350),
    .O(net_50320)
  );
  Odrv4 odrv_12_11_46351_50091 (
    .I(net_46351),
    .O(net_50091)
  );
  Odrv4 odrv_12_11_46352_50331 (
    .I(net_46352),
    .O(net_50331)
  );
  Odrv4 odrv_12_11_46353_50333 (
    .I(net_46353),
    .O(net_50333)
  );
  Odrv4 odrv_12_11_46354_50335 (
    .I(net_46354),
    .O(net_50335)
  );
  Odrv4 odrv_12_12_46474_50445 (
    .I(net_46474),
    .O(net_50445)
  );
  Odrv4 odrv_12_13_46596_39068 (
    .I(net_46596),
    .O(net_39068)
  );
  Odrv4 odrv_12_13_46596_46503 (
    .I(net_46596),
    .O(net_46503)
  );
  Odrv4 odrv_12_13_46596_46740 (
    .I(net_46596),
    .O(net_46740)
  );
  Odrv4 odrv_12_13_46596_46741 (
    .I(net_46596),
    .O(net_46741)
  );
  Odrv4 odrv_12_13_46596_50207 (
    .I(net_46596),
    .O(net_50207)
  );
  Odrv4 odrv_12_13_46596_50573 (
    .I(net_46596),
    .O(net_50573)
  );
  Odrv4 odrv_12_13_46599_50579 (
    .I(net_46599),
    .O(net_50579)
  );
  Odrv4 odrv_12_14_46717_46496 (
    .I(net_46717),
    .O(net_46496)
  );
  Odrv4 odrv_12_14_46723_50450 (
    .I(net_46723),
    .O(net_50450)
  );
  Odrv4 odrv_12_15_46840_50806 (
    .I(net_46840),
    .O(net_50806)
  );
  Odrv4 odrv_12_15_46841_43146 (
    .I(net_46841),
    .O(net_43146)
  );
  Odrv4 odrv_12_15_46841_46621 (
    .I(net_46841),
    .O(net_46621)
  );
  Odrv4 odrv_12_15_46841_46747 (
    .I(net_46841),
    .O(net_46747)
  );
  Odrv4 odrv_12_15_46841_46875 (
    .I(net_46841),
    .O(net_46875)
  );
  Odrv4 odrv_12_15_46841_50451 (
    .I(net_46841),
    .O(net_50451)
  );
  Odrv4 odrv_12_15_46842_39314 (
    .I(net_46842),
    .O(net_39314)
  );
  Odrv4 odrv_12_15_46842_46749 (
    .I(net_46842),
    .O(net_46749)
  );
  Odrv4 odrv_12_15_46842_46986 (
    .I(net_46842),
    .O(net_46986)
  );
  Odrv4 odrv_12_15_46842_50453 (
    .I(net_46842),
    .O(net_50453)
  );
  Odrv4 odrv_12_15_46842_50581 (
    .I(net_46842),
    .O(net_50581)
  );
  Odrv4 odrv_12_15_46842_50812 (
    .I(net_46842),
    .O(net_50812)
  );
  Odrv4 odrv_12_15_46843_39318 (
    .I(net_46843),
    .O(net_39318)
  );
  Odrv4 odrv_12_15_46843_46978 (
    .I(net_46843),
    .O(net_46978)
  );
  Odrv4 odrv_12_15_46843_50455 (
    .I(net_46843),
    .O(net_50455)
  );
  Odrv4 odrv_12_15_46843_50583 (
    .I(net_46843),
    .O(net_50583)
  );
  Odrv4 odrv_12_15_46847_43152 (
    .I(net_46847),
    .O(net_43152)
  );
  Odrv4 odrv_12_15_46847_46743 (
    .I(net_46847),
    .O(net_46743)
  );
  Odrv4 odrv_12_15_46847_46997 (
    .I(net_46847),
    .O(net_46997)
  );
  Odrv4 odrv_12_15_46847_50575 (
    .I(net_46847),
    .O(net_50575)
  );
  Odrv4 odrv_12_15_46847_50701 (
    .I(net_46847),
    .O(net_50701)
  );
  Odrv12 odrv_12_16_46965_49698 (
    .I(net_46965),
    .O(net_49698)
  );
  Odrv4 odrv_12_17_47092_46987 (
    .I(net_47092),
    .O(net_46987)
  );
  Odrv4 odrv_12_17_47093_46989 (
    .I(net_47093),
    .O(net_46989)
  );
  Odrv4 odrv_12_17_47093_50821 (
    .I(net_47093),
    .O(net_50821)
  );
  Odrv4 odrv_12_1_45078_45257 (
    .I(net_45078),
    .O(net_45257)
  );
  Odrv4 odrv_12_1_45078_49071 (
    .I(net_45078),
    .O(net_49071)
  );
  Odrv4 odrv_12_1_45078_49089 (
    .I(net_45078),
    .O(net_49089)
  );
  Odrv4 odrv_12_1_45079_49074 (
    .I(net_45079),
    .O(net_49074)
  );
  Odrv4 odrv_12_1_45079_49091 (
    .I(net_45079),
    .O(net_49091)
  );
  Odrv4 odrv_12_1_45080_49076 (
    .I(net_45080),
    .O(net_49076)
  );
  Odrv4 odrv_12_1_45080_49093 (
    .I(net_45080),
    .O(net_49093)
  );
  Odrv4 odrv_12_1_45081_49078 (
    .I(net_45081),
    .O(net_49078)
  );
  Odrv4 odrv_12_1_45081_49096 (
    .I(net_45081),
    .O(net_49096)
  );
  Odrv4 odrv_12_2_45206_45271 (
    .I(net_45206),
    .O(net_45271)
  );
  Odrv4 odrv_12_2_45206_49211 (
    .I(net_45206),
    .O(net_49211)
  );
  Odrv4 odrv_12_2_45208_37719 (
    .I(net_45208),
    .O(net_37719)
  );
  Odrv4 odrv_12_2_45208_45258 (
    .I(net_45208),
    .O(net_45258)
  );
  Odrv4 odrv_12_2_45208_45390 (
    .I(net_45208),
    .O(net_45390)
  );
  Odrv4 odrv_12_2_45209_45392 (
    .I(net_45209),
    .O(net_45392)
  );
  Odrv4 odrv_12_2_45209_49090 (
    .I(net_45209),
    .O(net_49090)
  );
  Odrv4 odrv_12_2_45209_49224 (
    .I(net_45209),
    .O(net_49224)
  );
  Odrv4 odrv_12_31_48810_48880 (
    .I(net_48810),
    .O(net_48880)
  );
  Odrv4 odrv_12_3_45368_37844 (
    .I(net_45368),
    .O(net_37844)
  );
  Odrv4 odrv_12_3_45368_41668 (
    .I(net_45368),
    .O(net_41668)
  );
  Odrv4 odrv_12_3_45368_45389 (
    .I(net_45368),
    .O(net_45389)
  );
  Odrv4 odrv_12_3_45368_45515 (
    .I(net_45368),
    .O(net_45515)
  );
  Odrv4 odrv_12_3_45368_49219 (
    .I(net_45368),
    .O(net_49219)
  );
  Odrv4 odrv_12_3_45368_49340 (
    .I(net_45368),
    .O(net_49340)
  );
  Odrv4 odrv_12_3_45370_41674 (
    .I(net_45370),
    .O(net_41674)
  );
  Odrv4 odrv_12_3_45370_45259 (
    .I(net_45370),
    .O(net_45259)
  );
  Odrv4 odrv_12_3_45370_49351 (
    .I(net_45370),
    .O(net_49351)
  );
  Odrv4 odrv_12_3_45371_45395 (
    .I(net_45371),
    .O(net_45395)
  );
  Odrv12 odrv_12_3_45371_48926 (
    .I(net_45371),
    .O(net_48926)
  );
  Odrv4 odrv_12_4_45488_45631 (
    .I(net_45488),
    .O(net_45631)
  );
  Odrv4 odrv_12_4_45489_45634 (
    .I(net_45489),
    .O(net_45634)
  );
  Odrv4 odrv_12_4_45493_49346 (
    .I(net_45493),
    .O(net_49346)
  );
  Odrv4 odrv_12_4_45494_45627 (
    .I(net_45494),
    .O(net_45627)
  );
  Odrv4 odrv_12_5_45610_49576 (
    .I(net_45610),
    .O(net_49576)
  );
  Odrv4 odrv_12_5_45612_45757 (
    .I(net_45612),
    .O(net_45757)
  );
  Odrv4 odrv_12_5_45615_49578 (
    .I(net_45615),
    .O(net_49578)
  );
  Odrv4 odrv_12_5_45616_49343 (
    .I(net_45616),
    .O(net_49343)
  );
  Odrv4 odrv_12_6_45737_38213 (
    .I(net_45737),
    .O(net_38213)
  );
  Odrv4 odrv_12_6_45737_45884 (
    .I(net_45737),
    .O(net_45884)
  );
  Odrv4 odrv_12_6_45738_45886 (
    .I(net_45738),
    .O(net_45886)
  );
  Odrv4 odrv_12_6_45739_45888 (
    .I(net_45739),
    .O(net_45888)
  );
  Odrv12 odrv_12_6_45739_48932 (
    .I(net_45739),
    .O(net_48932)
  );
  Odrv4 odrv_12_7_45859_45994 (
    .I(net_45859),
    .O(net_45994)
  );
  Odrv4 odrv_12_7_45860_42160 (
    .I(net_45860),
    .O(net_42160)
  );
  Odrv4 odrv_12_8_45979_49945 (
    .I(net_45979),
    .O(net_49945)
  );
  Odrv4 odrv_12_8_45983_49955 (
    .I(net_45983),
    .O(net_49955)
  );
  Odrv4 odrv_12_8_45984_49836 (
    .I(net_45984),
    .O(net_49836)
  );
  Odrv4 odrv_12_8_45986_46136 (
    .I(net_45986),
    .O(net_46136)
  );
  Odrv4 odrv_12_9_46102_42416 (
    .I(net_46102),
    .O(net_42416)
  );
  Odrv4 odrv_12_9_46107_50087 (
    .I(net_46107),
    .O(net_50087)
  );
  Odrv4 odrv_12_9_46108_42412 (
    .I(net_46108),
    .O(net_42412)
  );
  Odrv4 odrv_13_0_49034_49073 (
    .I(net_49034),
    .O(net_49073)
  );
  Odrv4 odrv_13_0_49034_49094 (
    .I(net_49034),
    .O(net_49094)
  );
  Odrv12 odrv_13_10_50056_53529 (
    .I(net_50056),
    .O(net_53529)
  );
  Odrv4 odrv_13_10_50060_53911 (
    .I(net_50060),
    .O(net_53911)
  );
  Odrv12 odrv_13_11_50180_53774 (
    .I(net_50180),
    .O(net_53774)
  );
  Odrv12 odrv_13_11_50181_53898 (
    .I(net_50181),
    .O(net_53898)
  );
  Odrv4 odrv_13_11_50183_54155 (
    .I(net_50183),
    .O(net_54155)
  );
  Odrv4 odrv_13_11_50184_49968 (
    .I(net_50184),
    .O(net_49968)
  );
  Odrv4 odrv_13_11_50185_50334 (
    .I(net_50185),
    .O(net_50334)
  );
  Odrv4 odrv_13_12_50303_46608 (
    .I(net_50303),
    .O(net_46608)
  );
  Odrv4 odrv_13_12_50309_54163 (
    .I(net_50309),
    .O(net_54163)
  );
  Odrv4 odrv_13_13_50426_50460 (
    .I(net_50426),
    .O(net_50460)
  );
  Odrv4 odrv_13_13_50429_54408 (
    .I(net_50429),
    .O(net_54408)
  );
  Odrv4 odrv_13_13_50431_50580 (
    .I(net_50431),
    .O(net_50580)
  );
  Odrv4 odrv_13_13_50432_54286 (
    .I(net_50432),
    .O(net_54286)
  );
  Odrv4 odrv_13_14_50548_50327 (
    .I(net_50548),
    .O(net_50327)
  );
  Odrv4 odrv_13_14_50549_46854 (
    .I(net_50549),
    .O(net_46854)
  );
  Odrv4 odrv_13_14_50549_50692 (
    .I(net_50549),
    .O(net_50692)
  );
  Odrv4 odrv_13_14_50549_54159 (
    .I(net_50549),
    .O(net_54159)
  );
  Odrv4 odrv_13_14_50549_54413 (
    .I(net_50549),
    .O(net_54413)
  );
  Odrv4 odrv_13_14_50549_54518 (
    .I(net_50549),
    .O(net_54518)
  );
  Odrv4 odrv_13_14_50551_50697 (
    .I(net_50551),
    .O(net_50697)
  );
  Odrv4 odrv_13_14_50552_43028 (
    .I(net_50552),
    .O(net_43028)
  );
  Odrv12 odrv_13_14_50553_53651 (
    .I(net_50553),
    .O(net_53651)
  );
  Odrv4 odrv_13_14_50554_46858 (
    .I(net_50554),
    .O(net_46858)
  );
  Odrv12 odrv_13_14_50555_53897 (
    .I(net_50555),
    .O(net_53897)
  );
  Odrv12 odrv_13_15_50671_54144 (
    .I(net_50671),
    .O(net_54144)
  );
  Odrv4 odrv_13_15_50672_50578 (
    .I(net_50672),
    .O(net_50578)
  );
  Odrv4 odrv_13_15_50675_54654 (
    .I(net_50675),
    .O(net_54654)
  );
  Odrv4 odrv_13_15_50676_54656 (
    .I(net_50676),
    .O(net_54656)
  );
  Odrv4 odrv_13_15_50677_54658 (
    .I(net_50677),
    .O(net_54658)
  );
  Odrv4 odrv_13_15_50678_50828 (
    .I(net_50678),
    .O(net_50828)
  );
  Odrv4 odrv_13_16_50797_43272 (
    .I(net_50797),
    .O(net_43272)
  );
  Odrv4 odrv_13_16_50797_50932 (
    .I(net_50797),
    .O(net_50932)
  );
  Odrv4 odrv_13_16_50797_50943 (
    .I(net_50797),
    .O(net_50943)
  );
  Odrv4 odrv_13_16_50797_54409 (
    .I(net_50797),
    .O(net_54409)
  );
  Odrv4 odrv_13_16_50797_54775 (
    .I(net_50797),
    .O(net_54775)
  );
  Odrv4 odrv_13_16_50798_54411 (
    .I(net_50798),
    .O(net_54411)
  );
  Odrv4 odrv_13_17_50924_43393 (
    .I(net_50924),
    .O(net_43393)
  );
  Odrv4 odrv_13_17_50924_47229 (
    .I(net_50924),
    .O(net_47229)
  );
  Odrv4 odrv_13_17_50924_50820 (
    .I(net_50924),
    .O(net_50820)
  );
  Odrv4 odrv_13_17_50924_50948 (
    .I(net_50924),
    .O(net_50948)
  );
  Odrv4 odrv_13_17_50924_51057 (
    .I(net_50924),
    .O(net_51057)
  );
  Odrv4 odrv_13_17_50924_54652 (
    .I(net_50924),
    .O(net_54652)
  );
  Odrv4 odrv_13_18_51040_51073 (
    .I(net_51040),
    .O(net_51073)
  );
  Odrv4 odrv_13_18_51043_43518 (
    .I(net_51043),
    .O(net_43518)
  );
  Odrv4 odrv_13_18_51045_51067 (
    .I(net_51045),
    .O(net_51067)
  );
  Odrv4 odrv_13_18_51047_51180 (
    .I(net_51047),
    .O(net_51180)
  );
  Odrv4 odrv_13_19_51170_51066 (
    .I(net_51170),
    .O(net_51066)
  );
  Odrv4 odrv_13_1_48911_49051 (
    .I(net_48911),
    .O(net_49051)
  );
  Odrv4 odrv_13_1_48911_49092 (
    .I(net_48911),
    .O(net_49092)
  );
  Odrv12 odrv_13_1_48911_52762 (
    .I(net_48911),
    .O(net_52762)
  );
  Odrv4 odrv_13_1_48914_41397 (
    .I(net_48914),
    .O(net_41397)
  );
  Odrv4 odrv_13_2_49038_53051 (
    .I(net_49038),
    .O(net_53051)
  );
  Odrv4 odrv_13_2_49040_52921 (
    .I(net_49040),
    .O(net_52921)
  );
  Odrv4 odrv_13_3_49196_49230 (
    .I(net_49196),
    .O(net_49230)
  );
  Odrv4 odrv_13_3_49196_53060 (
    .I(net_49196),
    .O(net_53060)
  );
  Odrv4 odrv_13_3_49196_53165 (
    .I(net_49196),
    .O(net_53165)
  );
  Odrv4 odrv_13_3_49200_53163 (
    .I(net_49200),
    .O(net_53163)
  );
  Odrv4 odrv_13_4_49318_49460 (
    .I(net_49318),
    .O(net_49460)
  );
  Odrv4 odrv_13_4_49319_53183 (
    .I(net_49319),
    .O(net_53183)
  );
  Odrv4 odrv_13_4_49320_41792 (
    .I(net_49320),
    .O(net_41792)
  );
  Odrv4 odrv_13_4_49320_49464 (
    .I(net_49320),
    .O(net_49464)
  );
  Odrv4 odrv_13_4_49320_53290 (
    .I(net_49320),
    .O(net_53290)
  );
  Odrv4 odrv_13_4_49321_41796 (
    .I(net_49321),
    .O(net_41796)
  );
  Odrv4 odrv_13_4_49321_49456 (
    .I(net_49321),
    .O(net_49456)
  );
  Odrv4 odrv_13_4_49321_49467 (
    .I(net_49321),
    .O(net_49467)
  );
  Odrv4 odrv_13_4_49322_49469 (
    .I(net_49322),
    .O(net_49469)
  );
  Odrv4 odrv_13_4_49322_53294 (
    .I(net_49322),
    .O(net_53294)
  );
  Odrv4 odrv_13_4_49322_53301 (
    .I(net_49322),
    .O(net_53301)
  );
  Odrv4 odrv_13_4_49325_53053 (
    .I(net_49325),
    .O(net_53053)
  );
  Odrv4 odrv_13_5_49446_49468 (
    .I(net_49446),
    .O(net_49468)
  );
  Odrv4 odrv_13_5_49447_53428 (
    .I(net_49447),
    .O(net_53428)
  );
  Odrv4 odrv_13_6_49564_53530 (
    .I(net_49564),
    .O(net_53530)
  );
  Odrv4 odrv_13_6_49565_53534 (
    .I(net_49565),
    .O(net_53534)
  );
  Odrv4 odrv_13_6_49566_49710 (
    .I(net_49566),
    .O(net_49710)
  );
  Odrv4 odrv_13_6_49567_53179 (
    .I(net_49567),
    .O(net_53179)
  );
  Odrv4 odrv_13_6_49568_53540 (
    .I(net_49568),
    .O(net_53540)
  );
  Odrv4 odrv_13_6_49569_53532 (
    .I(net_49569),
    .O(net_53532)
  );
  Odrv4 odrv_13_6_49570_42048 (
    .I(net_49570),
    .O(net_42048)
  );
  Odrv4 odrv_13_6_49571_45876 (
    .I(net_49571),
    .O(net_45876)
  );
  Odrv4 odrv_13_7_49688_53657 (
    .I(net_49688),
    .O(net_53657)
  );
  Odrv4 odrv_13_7_49689_53666 (
    .I(net_49689),
    .O(net_53666)
  );
  Odrv4 odrv_13_7_49691_53670 (
    .I(net_49691),
    .O(net_53670)
  );
  Odrv4 odrv_13_7_49692_53672 (
    .I(net_49692),
    .O(net_53672)
  );
  Odrv4 odrv_13_7_49694_49827 (
    .I(net_49694),
    .O(net_49827)
  );
  Odrv4 odrv_13_8_49810_46124 (
    .I(net_49810),
    .O(net_46124)
  );
  Odrv4 odrv_13_8_49811_53780 (
    .I(net_49811),
    .O(net_53780)
  );
  Odrv4 odrv_13_8_49812_49956 (
    .I(net_49812),
    .O(net_49956)
  );
  Odrv4 odrv_13_8_49814_46114 (
    .I(net_49814),
    .O(net_46114)
  );
  Odrv4 odrv_13_8_49817_49841 (
    .I(net_49817),
    .O(net_49841)
  );
  Odrv4 odrv_14_10_53887_54029 (
    .I(net_53887),
    .O(net_54029)
  );
  Odrv4 odrv_14_10_53888_54031 (
    .I(net_53888),
    .O(net_54031)
  );
  Odrv4 odrv_14_10_53888_57751 (
    .I(net_53888),
    .O(net_57751)
  );
  Odrv4 odrv_14_10_53889_54033 (
    .I(net_53889),
    .O(net_54033)
  );
  Odrv4 odrv_14_10_53890_54025 (
    .I(net_53890),
    .O(net_54025)
  );
  Odrv4 odrv_14_10_53891_53674 (
    .I(net_53891),
    .O(net_53674)
  );
  Odrv12 odrv_14_10_53892_54019 (
    .I(net_53892),
    .O(net_54019)
  );
  Odrv4 odrv_14_10_53892_57743 (
    .I(net_53892),
    .O(net_57743)
  );
  Odrv4 odrv_14_10_53893_57619 (
    .I(net_53893),
    .O(net_57619)
  );
  Odrv4 odrv_14_10_53893_57745 (
    .I(net_53893),
    .O(net_57745)
  );
  Odrv4 odrv_14_10_53894_54027 (
    .I(net_53894),
    .O(net_54027)
  );
  Odrv4 odrv_14_10_53894_57747 (
    .I(net_53894),
    .O(net_57747)
  );
  Odrv4 odrv_14_11_54010_57746 (
    .I(net_54010),
    .O(net_57746)
  );
  Odrv4 odrv_14_11_54013_57752 (
    .I(net_54013),
    .O(net_57752)
  );
  Odrv4 odrv_14_11_54014_50314 (
    .I(net_54014),
    .O(net_50314)
  );
  Odrv4 odrv_14_11_54017_57744 (
    .I(net_54017),
    .O(net_57744)
  );
  Odrv4 odrv_14_12_54137_53920 (
    .I(net_54137),
    .O(net_53920)
  );
  Odrv4 odrv_14_12_54137_54284 (
    .I(net_54137),
    .O(net_54284)
  );
  Odrv4 odrv_14_13_54256_58221 (
    .I(net_54256),
    .O(net_58221)
  );
  Odrv12 odrv_14_13_54258_35232 (
    .I(net_54258),
    .O(net_35232)
  );
  Odrv4 odrv_14_13_54258_46730 (
    .I(net_54258),
    .O(net_46730)
  );
  Odrv4 odrv_14_13_54258_57996 (
    .I(net_54258),
    .O(net_57996)
  );
  Odrv4 odrv_14_13_54259_58236 (
    .I(net_54259),
    .O(net_58236)
  );
  Odrv4 odrv_14_13_54261_58223 (
    .I(net_54261),
    .O(net_58223)
  );
  Odrv12 odrv_14_13_54262_57482 (
    .I(net_54262),
    .O(net_57482)
  );
  Odrv4 odrv_14_13_54262_58114 (
    .I(net_54262),
    .O(net_58114)
  );
  Odrv4 odrv_14_13_54263_46732 (
    .I(net_54263),
    .O(net_46732)
  );
  Odrv4 odrv_14_13_54263_54396 (
    .I(net_54263),
    .O(net_54396)
  );
  Odrv4 odrv_14_13_54263_58116 (
    .I(net_54263),
    .O(net_58116)
  );
  Odrv4 odrv_14_14_54379_57987 (
    .I(net_54379),
    .O(net_57987)
  );
  Odrv4 odrv_14_14_54379_58241 (
    .I(net_54379),
    .O(net_58241)
  );
  Odrv4 odrv_14_14_54381_58350 (
    .I(net_54381),
    .O(net_58350)
  );
  Odrv4 odrv_14_14_54381_58357 (
    .I(net_54381),
    .O(net_58357)
  );
  Odrv4 odrv_14_14_54383_58354 (
    .I(net_54383),
    .O(net_58354)
  );
  Odrv4 odrv_14_14_54383_58361 (
    .I(net_54383),
    .O(net_58361)
  );
  Odrv4 odrv_14_14_54384_58346 (
    .I(net_54384),
    .O(net_58346)
  );
  Odrv4 odrv_14_14_54384_58363 (
    .I(net_54384),
    .O(net_58363)
  );
  Odrv12 odrv_14_14_54385_57605 (
    .I(net_54385),
    .O(net_57605)
  );
  Odrv4 odrv_14_14_54386_50691 (
    .I(net_54386),
    .O(net_50691)
  );
  Odrv4 odrv_14_14_54386_58367 (
    .I(net_54386),
    .O(net_58367)
  );
  Odrv12 odrv_14_15_54503_58096 (
    .I(net_54503),
    .O(net_58096)
  );
  Odrv4 odrv_14_15_54504_46976 (
    .I(net_54504),
    .O(net_46976)
  );
  Odrv4 odrv_14_15_54506_54289 (
    .I(net_54506),
    .O(net_54289)
  );
  Odrv4 odrv_14_16_54627_58596 (
    .I(net_54627),
    .O(net_58596)
  );
  Odrv4 odrv_14_16_54628_58605 (
    .I(net_54628),
    .O(net_58605)
  );
  Odrv4 odrv_14_16_54629_50929 (
    .I(net_54629),
    .O(net_50929)
  );
  Odrv4 odrv_14_16_54630_58243 (
    .I(net_54630),
    .O(net_58243)
  );
  Odrv4 odrv_14_16_54631_54780 (
    .I(net_54631),
    .O(net_54780)
  );
  Odrv4 odrv_14_16_54632_54765 (
    .I(net_54632),
    .O(net_54765)
  );
  Odrv4 odrv_14_17_54748_58713 (
    .I(net_54748),
    .O(net_58713)
  );
  Odrv4 odrv_14_17_54749_58358 (
    .I(net_54749),
    .O(net_58358)
  );
  Odrv4 odrv_14_17_54749_58486 (
    .I(net_54749),
    .O(net_58486)
  );
  Odrv4 odrv_14_17_54749_58717 (
    .I(net_54749),
    .O(net_58717)
  );
  Odrv4 odrv_14_18_54872_58481 (
    .I(net_54872),
    .O(net_58481)
  );
  Odrv4 odrv_14_18_54873_58483 (
    .I(net_54873),
    .O(net_58483)
  );
  Odrv4 odrv_14_18_54876_54660 (
    .I(net_54876),
    .O(net_54660)
  );
  Odrv4 odrv_14_18_54876_58489 (
    .I(net_54876),
    .O(net_58489)
  );
  Odrv4 odrv_14_18_54877_54772 (
    .I(net_54877),
    .O(net_54772)
  );
  Odrv4 odrv_14_18_54877_58603 (
    .I(net_54877),
    .O(net_58603)
  );
  Odrv4 odrv_14_19_54997_54905 (
    .I(net_54997),
    .O(net_54905)
  );
  Odrv4 odrv_14_1_52745_45228 (
    .I(net_52745),
    .O(net_45228)
  );
  Odrv4 odrv_14_2_52870_56883 (
    .I(net_52870),
    .O(net_56883)
  );
  Odrv4 odrv_14_4_53151_45623 (
    .I(net_53151),
    .O(net_45623)
  );
  Odrv4 odrv_14_4_53151_53295 (
    .I(net_53151),
    .O(net_53295)
  );
  Odrv4 odrv_14_4_53151_53296 (
    .I(net_53151),
    .O(net_53296)
  );
  Odrv4 odrv_14_4_53151_56889 (
    .I(net_53151),
    .O(net_56889)
  );
  Odrv4 odrv_14_4_53153_57003 (
    .I(net_53153),
    .O(net_57003)
  );
  Odrv4 odrv_14_4_53155_57135 (
    .I(net_53155),
    .O(net_57135)
  );
  Odrv4 odrv_14_4_53156_49461 (
    .I(net_53156),
    .O(net_49461)
  );
  Odrv4 odrv_14_5_53272_57008 (
    .I(net_53272),
    .O(net_57008)
  );
  Odrv4 odrv_14_6_53396_57364 (
    .I(net_53396),
    .O(net_57364)
  );
  Odrv12 odrv_14_6_53399_57356 (
    .I(net_53399),
    .O(net_57356)
  );
  Odrv4 odrv_14_6_53399_57370 (
    .I(net_53399),
    .O(net_57370)
  );
  Odrv4 odrv_14_6_53401_45879 (
    .I(net_53401),
    .O(net_45879)
  );
  Odrv4 odrv_14_7_53521_45996 (
    .I(net_53521),
    .O(net_45996)
  );
  Odrv4 odrv_14_7_53524_49828 (
    .I(net_53524),
    .O(net_49828)
  );
  Odrv4 odrv_14_7_53524_53654 (
    .I(net_53524),
    .O(net_53654)
  );
  Odrv4 odrv_14_7_53524_53673 (
    .I(net_53524),
    .O(net_53673)
  );
  Odrv4 odrv_14_8_53641_57606 (
    .I(net_53641),
    .O(net_57606)
  );
  Odrv4 odrv_14_8_53642_57610 (
    .I(net_53642),
    .O(net_57610)
  );
  Odrv4 odrv_14_8_53643_53550 (
    .I(net_53643),
    .O(net_53550)
  );
  Odrv4 odrv_14_8_53643_53788 (
    .I(net_53643),
    .O(net_53788)
  );
  Odrv4 odrv_14_8_53644_46119 (
    .I(net_53644),
    .O(net_46119)
  );
  Odrv4 odrv_14_8_53644_53552 (
    .I(net_53644),
    .O(net_53552)
  );
  Odrv4 odrv_14_8_53644_53779 (
    .I(net_53644),
    .O(net_53779)
  );
  Odrv4 odrv_14_8_53644_57621 (
    .I(net_53644),
    .O(net_57621)
  );
  Odrv4 odrv_14_8_53645_46121 (
    .I(net_53645),
    .O(net_46121)
  );
  Odrv4 odrv_14_8_53647_53777 (
    .I(net_53647),
    .O(net_53777)
  );
  Odrv4 odrv_14_8_53648_46117 (
    .I(net_53648),
    .O(net_46117)
  );
  Odrv4 odrv_14_8_53648_53798 (
    .I(net_53648),
    .O(net_53798)
  );
  Odrv4 odrv_14_8_53648_57629 (
    .I(net_53648),
    .O(net_57629)
  );
  Odrv4 odrv_14_9_53770_57750 (
    .I(net_53770),
    .O(net_57750)
  );
  Odrv4 odrv_15_0_56693_56738 (
    .I(net_56693),
    .O(net_56738)
  );
  Odrv4 odrv_15_10_57724_54030 (
    .I(net_57724),
    .O(net_54030)
  );
  Odrv4 odrv_15_11_57840_57982 (
    .I(net_57840),
    .O(net_57982)
  );
  Odrv4 odrv_15_11_57840_61702 (
    .I(net_57840),
    .O(net_61702)
  );
  Odrv4 odrv_15_11_57840_61805 (
    .I(net_57840),
    .O(net_61805)
  );
  Odrv4 odrv_15_11_57843_57978 (
    .I(net_57843),
    .O(net_57978)
  );
  Odrv4 odrv_15_11_57845_50323 (
    .I(net_57845),
    .O(net_50323)
  );
  Odrv4 odrv_15_11_57846_54151 (
    .I(net_57846),
    .O(net_54151)
  );
  Odrv4 odrv_15_11_57846_57741 (
    .I(net_57846),
    .O(net_57741)
  );
  Odrv4 odrv_15_11_57846_57995 (
    .I(net_57846),
    .O(net_57995)
  );
  Odrv4 odrv_15_11_57846_61826 (
    .I(net_57846),
    .O(net_61826)
  );
  Odrv4 odrv_15_12_57963_61825 (
    .I(net_57963),
    .O(net_61825)
  );
  Odrv4 odrv_15_12_57968_57990 (
    .I(net_57968),
    .O(net_57990)
  );
  Odrv4 odrv_15_13_58090_50567 (
    .I(net_58090),
    .O(net_50567)
  );
  Odrv4 odrv_15_13_58092_58115 (
    .I(net_58092),
    .O(net_58115)
  );
  Odrv4 odrv_15_14_58209_62174 (
    .I(net_58209),
    .O(net_62174)
  );
  Odrv4 odrv_15_14_58210_54516 (
    .I(net_58210),
    .O(net_54516)
  );
  Odrv4 odrv_15_14_58211_58355 (
    .I(net_58211),
    .O(net_58355)
  );
  Odrv4 odrv_15_14_58211_62180 (
    .I(net_58211),
    .O(net_62180)
  );
  Odrv4 odrv_15_14_58212_61823 (
    .I(net_58212),
    .O(net_61823)
  );
  Odrv4 odrv_15_14_58212_61951 (
    .I(net_58212),
    .O(net_61951)
  );
  Odrv4 odrv_15_14_58213_54514 (
    .I(net_58213),
    .O(net_54514)
  );
  Odrv4 odrv_15_14_58214_57998 (
    .I(net_58214),
    .O(net_57998)
  );
  Odrv4 odrv_15_14_58215_54520 (
    .I(net_58215),
    .O(net_54520)
  );
  Odrv4 odrv_15_14_58215_58110 (
    .I(net_58215),
    .O(net_58110)
  );
  Odrv4 odrv_15_14_58216_50686 (
    .I(net_58216),
    .O(net_50686)
  );
  Odrv4 odrv_15_14_58216_62197 (
    .I(net_58216),
    .O(net_62197)
  );
  Odrv4 odrv_15_15_58332_58365 (
    .I(net_58332),
    .O(net_58365)
  );
  Odrv4 odrv_15_15_58332_62068 (
    .I(net_58332),
    .O(net_62068)
  );
  Odrv4 odrv_15_15_58336_61948 (
    .I(net_58336),
    .O(net_61948)
  );
  Odrv4 odrv_15_15_58338_58233 (
    .I(net_58338),
    .O(net_58233)
  );
  Odrv4 odrv_15_15_58339_62066 (
    .I(net_58339),
    .O(net_62066)
  );
  Odrv4 odrv_15_16_58458_58604 (
    .I(net_58458),
    .O(net_58604)
  );
  Odrv4 odrv_15_16_58461_58610 (
    .I(net_58461),
    .O(net_58610)
  );
  Odrv4 odrv_15_17_58579_62547 (
    .I(net_58579),
    .O(net_62547)
  );
  Odrv4 odrv_15_18_58705_58488 (
    .I(net_58705),
    .O(net_58488)
  );
  Odrv4 odrv_15_2_56703_56757 (
    .I(net_56703),
    .O(net_56757)
  );
  Odrv4 odrv_15_3_56860_49337 (
    .I(net_56860),
    .O(net_49337)
  );
  Odrv4 odrv_15_4_56980_53286 (
    .I(net_56980),
    .O(net_53286)
  );
  Odrv4 odrv_15_4_56982_60952 (
    .I(net_56982),
    .O(net_60952)
  );
  Odrv4 odrv_15_4_56982_60959 (
    .I(net_56982),
    .O(net_60959)
  );
  Odrv4 odrv_15_4_56983_53284 (
    .I(net_56983),
    .O(net_53284)
  );
  Odrv4 odrv_15_4_56983_60961 (
    .I(net_56983),
    .O(net_60961)
  );
  Odrv4 odrv_15_4_56984_53288 (
    .I(net_56984),
    .O(net_53288)
  );
  Odrv4 odrv_15_4_56985_57134 (
    .I(net_56985),
    .O(net_57134)
  );
  Odrv4 odrv_15_4_56985_60837 (
    .I(net_56985),
    .O(net_60837)
  );
  Odrv4 odrv_15_5_57102_57007 (
    .I(net_57102),
    .O(net_57007)
  );
  Odrv4 odrv_15_5_57102_60964 (
    .I(net_57102),
    .O(net_60964)
  );
  Odrv4 odrv_15_5_57103_57009 (
    .I(net_57103),
    .O(net_57009)
  );
  Odrv4 odrv_15_5_57103_57137 (
    .I(net_57103),
    .O(net_57137)
  );
  Odrv12 odrv_15_5_57104_60411 (
    .I(net_57104),
    .O(net_60411)
  );
  Odrv4 odrv_15_5_57104_60842 (
    .I(net_57104),
    .O(net_60842)
  );
  Odrv4 odrv_15_5_57105_60844 (
    .I(net_57105),
    .O(net_60844)
  );
  Odrv4 odrv_15_5_57106_53407 (
    .I(net_57106),
    .O(net_53407)
  );
  Odrv4 odrv_15_5_57107_53411 (
    .I(net_57107),
    .O(net_53411)
  );
  Odrv4 odrv_15_5_57108_60834 (
    .I(net_57108),
    .O(net_60834)
  );
  Odrv4 odrv_15_5_57108_60960 (
    .I(net_57108),
    .O(net_60960)
  );
  Odrv4 odrv_15_5_57109_53415 (
    .I(net_57109),
    .O(net_53415)
  );
  Odrv4 odrv_15_6_57226_61194 (
    .I(net_57226),
    .O(net_61194)
  );
  Odrv4 odrv_15_6_57228_49704 (
    .I(net_57228),
    .O(net_49704)
  );
  Odrv4 odrv_15_6_57230_49708 (
    .I(net_57230),
    .O(net_49708)
  );
  Odrv4 odrv_15_6_57231_57126 (
    .I(net_57231),
    .O(net_57126)
  );
  Odrv4 odrv_15_8_57471_57250 (
    .I(net_57471),
    .O(net_57250)
  );
  Odrv4 odrv_15_8_57471_57504 (
    .I(net_57471),
    .O(net_57504)
  );
  Odrv4 odrv_15_8_57471_57613 (
    .I(net_57471),
    .O(net_57613)
  );
  Odrv4 odrv_15_8_57472_53778 (
    .I(net_57472),
    .O(net_53778)
  );
  Odrv4 odrv_15_8_57472_61081 (
    .I(net_57472),
    .O(net_61081)
  );
  Odrv4 odrv_15_8_57472_61335 (
    .I(net_57472),
    .O(net_61335)
  );
  Odrv4 odrv_15_8_57473_57618 (
    .I(net_57473),
    .O(net_57618)
  );
  Odrv4 odrv_15_8_57474_57609 (
    .I(net_57474),
    .O(net_57609)
  );
  Odrv4 odrv_15_8_57474_61213 (
    .I(net_57474),
    .O(net_61213)
  );
  Odrv4 odrv_15_8_57475_49952 (
    .I(net_57475),
    .O(net_49952)
  );
  Odrv4 odrv_15_8_57475_53776 (
    .I(net_57475),
    .O(net_53776)
  );
  Odrv4 odrv_15_9_57594_53909 (
    .I(net_57594),
    .O(net_53909)
  );
  Odrv4 odrv_15_9_57595_61204 (
    .I(net_57595),
    .O(net_61204)
  );
  Odrv4 odrv_15_9_57596_61572 (
    .I(net_57596),
    .O(net_61572)
  );
  Odrv4 odrv_15_9_57597_61574 (
    .I(net_57597),
    .O(net_61574)
  );
  Odrv4 odrv_15_9_57598_61576 (
    .I(net_57598),
    .O(net_61576)
  );
  Odrv4 odrv_15_9_57600_53905 (
    .I(net_57600),
    .O(net_53905)
  );
  Odrv4 odrv_16_10_61547_65284 (
    .I(net_61547),
    .O(net_65284)
  );
  Odrv4 odrv_16_10_61547_65410 (
    .I(net_61547),
    .O(net_65410)
  );
  Odrv4 odrv_16_10_61549_65288 (
    .I(net_61549),
    .O(net_65288)
  );
  Odrv4 odrv_16_10_61550_65290 (
    .I(net_61550),
    .O(net_65290)
  );
  Odrv4 odrv_16_10_61550_65528 (
    .I(net_61550),
    .O(net_65528)
  );
  Odrv4 odrv_16_10_61551_65530 (
    .I(net_61551),
    .O(net_65530)
  );
  Odrv4 odrv_16_10_61552_65532 (
    .I(net_61552),
    .O(net_65532)
  );
  Odrv4 odrv_16_10_61553_65406 (
    .I(net_61553),
    .O(net_65406)
  );
  Odrv4 odrv_16_10_61554_65408 (
    .I(net_61554),
    .O(net_65408)
  );
  Odrv12 odrv_16_11_61671_65265 (
    .I(net_61671),
    .O(net_65265)
  );
  Odrv4 odrv_16_11_61672_54146 (
    .I(net_61672),
    .O(net_54146)
  );
  Odrv4 odrv_16_11_61672_65411 (
    .I(net_61672),
    .O(net_65411)
  );
  Odrv12 odrv_16_11_61673_65511 (
    .I(net_61673),
    .O(net_65511)
  );
  Odrv4 odrv_16_11_61674_57975 (
    .I(net_61674),
    .O(net_57975)
  );
  Odrv4 odrv_16_11_61674_65646 (
    .I(net_61674),
    .O(net_65646)
  );
  Odrv4 odrv_16_11_61676_61571 (
    .I(net_61676),
    .O(net_61571)
  );
  Odrv4 odrv_16_11_61677_61573 (
    .I(net_61677),
    .O(net_61573)
  );
  Odrv4 odrv_16_12_61795_61939 (
    .I(net_61795),
    .O(net_61939)
  );
  Odrv4 odrv_16_12_61796_61578 (
    .I(net_61796),
    .O(net_61578)
  );
  Odrv4 odrv_16_12_61799_61929 (
    .I(net_61799),
    .O(net_61929)
  );
  Odrv4 odrv_16_12_61800_58106 (
    .I(net_61800),
    .O(net_58106)
  );
  Odrv4 odrv_16_13_61923_65651 (
    .I(net_61923),
    .O(net_65651)
  );
  Odrv4 odrv_16_13_61923_65777 (
    .I(net_61923),
    .O(net_65777)
  );
  Odrv4 odrv_16_15_62165_62073 (
    .I(net_62165),
    .O(net_62073)
  );
  Odrv4 odrv_16_15_62166_58467 (
    .I(net_62166),
    .O(net_58467)
  );
  Odrv4 odrv_16_15_62167_65781 (
    .I(net_62167),
    .O(net_65781)
  );
  Odrv4 odrv_16_15_62167_66130 (
    .I(net_62167),
    .O(net_66130)
  );
  Odrv4 odrv_16_15_62168_62298 (
    .I(net_62168),
    .O(net_62298)
  );
  Odrv4 odrv_16_16_62285_58600 (
    .I(net_62285),
    .O(net_58600)
  );
  Odrv4 odrv_16_16_62286_58592 (
    .I(net_62286),
    .O(net_58592)
  );
  Odrv4 odrv_16_16_62289_66261 (
    .I(net_62289),
    .O(net_66261)
  );
  Odrv4 odrv_16_16_62290_65904 (
    .I(net_62290),
    .O(net_65904)
  );
  Odrv4 odrv_16_16_62291_54771 (
    .I(net_62291),
    .O(net_54771)
  );
  Odrv4 odrv_16_17_62408_62187 (
    .I(net_62408),
    .O(net_62187)
  );
  Odrv4 odrv_16_17_62409_66019 (
    .I(net_62409),
    .O(net_66019)
  );
  Odrv4 odrv_16_17_62410_62555 (
    .I(net_62410),
    .O(net_62555)
  );
  Odrv4 odrv_16_17_62411_54888 (
    .I(net_62411),
    .O(net_54888)
  );
  Odrv4 odrv_16_17_62411_62193 (
    .I(net_62411),
    .O(net_62193)
  );
  Odrv4 odrv_16_17_62412_66025 (
    .I(net_62412),
    .O(net_66025)
  );
  Odrv4 odrv_16_17_62413_66393 (
    .I(net_62413),
    .O(net_66393)
  );
  Odrv4 odrv_16_17_62414_66141 (
    .I(net_62414),
    .O(net_66141)
  );
  Odrv4 odrv_16_17_62415_62548 (
    .I(net_62415),
    .O(net_62548)
  );
  Odrv12 odrv_16_18_62531_65020 (
    .I(net_62531),
    .O(net_65020)
  );
  Odrv4 odrv_16_2_60530_60701 (
    .I(net_60530),
    .O(net_60701)
  );
  Odrv4 odrv_16_3_60688_53162 (
    .I(net_60688),
    .O(net_53162)
  );
  Odrv4 odrv_16_3_60688_60590 (
    .I(net_60688),
    .O(net_60590)
  );
  Odrv4 odrv_16_3_60688_60833 (
    .I(net_60688),
    .O(net_60833)
  );
  Odrv12 odrv_16_3_60688_64260 (
    .I(net_60688),
    .O(net_64260)
  );
  Odrv4 odrv_16_3_60688_64658 (
    .I(net_60688),
    .O(net_64658)
  );
  Odrv4 odrv_16_3_60688_64665 (
    .I(net_60688),
    .O(net_64665)
  );
  Odrv4 odrv_16_3_60689_60835 (
    .I(net_60689),
    .O(net_60835)
  );
  Odrv4 odrv_16_3_60689_64424 (
    .I(net_60689),
    .O(net_64424)
  );
  Odrv4 odrv_16_3_60689_64660 (
    .I(net_60689),
    .O(net_64660)
  );
  Odrv4 odrv_16_4_60810_64674 (
    .I(net_60810),
    .O(net_64674)
  );
  Odrv4 odrv_16_4_60811_60956 (
    .I(net_60811),
    .O(net_60956)
  );
  Odrv4 odrv_16_4_60812_60958 (
    .I(net_60812),
    .O(net_60958)
  );
  Odrv4 odrv_16_4_60813_64792 (
    .I(net_60813),
    .O(net_64792)
  );
  Odrv4 odrv_16_4_60814_64666 (
    .I(net_60814),
    .O(net_64666)
  );
  Odrv4 odrv_16_4_60815_64796 (
    .I(net_60815),
    .O(net_64796)
  );
  Odrv4 odrv_16_4_60816_60966 (
    .I(net_60816),
    .O(net_60966)
  );
  Odrv4 odrv_16_5_60932_60965 (
    .I(net_60932),
    .O(net_60965)
  );
  Odrv4 odrv_16_5_60933_60967 (
    .I(net_60933),
    .O(net_60967)
  );
  Odrv4 odrv_16_5_60934_61079 (
    .I(net_60934),
    .O(net_61079)
  );
  Odrv4 odrv_16_5_60935_64913 (
    .I(net_60935),
    .O(net_64913)
  );
  Odrv4 odrv_16_5_60937_61085 (
    .I(net_60937),
    .O(net_61085)
  );
  Odrv4 odrv_16_6_61056_64920 (
    .I(net_61056),
    .O(net_64920)
  );
  Odrv4 odrv_16_6_61057_61201 (
    .I(net_61057),
    .O(net_61201)
  );
  Odrv4 odrv_16_6_61058_64798 (
    .I(net_61058),
    .O(net_64798)
  );
  Odrv4 odrv_16_6_61059_57360 (
    .I(net_61059),
    .O(net_57360)
  );
  Odrv4 odrv_16_6_61060_61208 (
    .I(net_61060),
    .O(net_61208)
  );
  Odrv4 odrv_16_6_61061_57366 (
    .I(net_61061),
    .O(net_57366)
  );
  Odrv4 odrv_16_6_61062_61212 (
    .I(net_61062),
    .O(net_61212)
  );
  Odrv4 odrv_16_7_61178_65144 (
    .I(net_61178),
    .O(net_65144)
  );
  Odrv4 odrv_16_7_61179_65148 (
    .I(net_61179),
    .O(net_65148)
  );
  Odrv4 odrv_16_7_61180_61324 (
    .I(net_61180),
    .O(net_61324)
  );
  Odrv4 odrv_16_7_61181_61316 (
    .I(net_61181),
    .O(net_61316)
  );
  Odrv4 odrv_16_7_61183_61205 (
    .I(net_61183),
    .O(net_61205)
  );
  Odrv4 odrv_16_7_61184_64911 (
    .I(net_61184),
    .O(net_64911)
  );
  Odrv4 odrv_16_7_61184_65037 (
    .I(net_61184),
    .O(net_65037)
  );
  Odrv4 odrv_16_7_61184_65165 (
    .I(net_61184),
    .O(net_65165)
  );
  Odrv4 odrv_16_7_61185_57491 (
    .I(net_61185),
    .O(net_57491)
  );
  Odrv4 odrv_16_8_61302_61336 (
    .I(net_61302),
    .O(net_61336)
  );
  Odrv4 odrv_16_8_61305_61452 (
    .I(net_61305),
    .O(net_61452)
  );
  Odrv4 odrv_16_9_61425_57731 (
    .I(net_61425),
    .O(net_57731)
  );
  Odrv4 odrv_16_9_61425_61459 (
    .I(net_61425),
    .O(net_61459)
  );
  Odrv12 odrv_16_9_61426_42402 (
    .I(net_61426),
    .O(net_42402)
  );
  Odrv4 odrv_16_9_61428_57729 (
    .I(net_61428),
    .O(net_57729)
  );
  Odrv4 odrv_16_9_61428_65279 (
    .I(net_61428),
    .O(net_65279)
  );
  Odrv4 odrv_16_9_61429_53908 (
    .I(net_61429),
    .O(net_53908)
  );
  Odrv4 odrv_16_9_61429_61577 (
    .I(net_61429),
    .O(net_61577)
  );
  Odrv4 odrv_16_9_61430_61325 (
    .I(net_61430),
    .O(net_61325)
  );
  Odrv4 odrv_16_9_61431_53902 (
    .I(net_61431),
    .O(net_53902)
  );
  Odrv4 odrv_17_0_64354_56601 (
    .I(net_64354),
    .O(net_56601)
  );
  Odrv4 odrv_17_0_64354_64408 (
    .I(net_64354),
    .O(net_64408)
  );
  Odrv12 odrv_17_10_65381_42526 (
    .I(net_65381),
    .O(net_42526)
  );
  Odrv4 odrv_17_10_65382_61682 (
    .I(net_65382),
    .O(net_61682)
  );
  Odrv4 odrv_17_10_65383_61686 (
    .I(net_65383),
    .O(net_61686)
  );
  Odrv4 odrv_17_10_65383_65167 (
    .I(net_65383),
    .O(net_65167)
  );
  Odrv4 odrv_17_10_65383_65405 (
    .I(net_65383),
    .O(net_65405)
  );
  Odrv4 odrv_17_10_65383_68997 (
    .I(net_65383),
    .O(net_68997)
  );
  Odrv4 odrv_17_11_65507_65402 (
    .I(net_65507),
    .O(net_65402)
  );
  Odrv12 odrv_17_11_65508_68850 (
    .I(net_65508),
    .O(net_68850)
  );
  Odrv4 odrv_17_13_65748_69717 (
    .I(net_65748),
    .O(net_69717)
  );
  Odrv4 odrv_17_14_65870_69836 (
    .I(net_65870),
    .O(net_69836)
  );
  Odrv4 odrv_17_14_65874_66021 (
    .I(net_65874),
    .O(net_66021)
  );
  Odrv4 odrv_17_15_65994_69604 (
    .I(net_65994),
    .O(net_69604)
  );
  Odrv4 odrv_17_15_65995_69965 (
    .I(net_65995),
    .O(net_69965)
  );
  Odrv4 odrv_17_15_65997_69610 (
    .I(net_65997),
    .O(net_69610)
  );
  Odrv4 odrv_17_15_65999_65894 (
    .I(net_65999),
    .O(net_65894)
  );
  Odrv4 odrv_17_16_66118_65899 (
    .I(net_66118),
    .O(net_65899)
  );
  Odrv4 odrv_17_16_66119_65901 (
    .I(net_66119),
    .O(net_65901)
  );
  Odrv4 odrv_17_16_66120_65903 (
    .I(net_66120),
    .O(net_65903)
  );
  Odrv4 odrv_17_16_66121_65905 (
    .I(net_66121),
    .O(net_65905)
  );
  Odrv4 odrv_17_16_66122_66017 (
    .I(net_66122),
    .O(net_66017)
  );
  Odrv4 odrv_17_17_66240_69850 (
    .I(net_66240),
    .O(net_69850)
  );
  Odrv4 odrv_17_17_66243_58720 (
    .I(net_66243),
    .O(net_58720)
  );
  Odrv4 odrv_17_17_66243_62543 (
    .I(net_66243),
    .O(net_62543)
  );
  Odrv4 odrv_17_17_66245_69972 (
    .I(net_66245),
    .O(net_69972)
  );
  Odrv4 odrv_17_17_66246_58716 (
    .I(net_66246),
    .O(net_58716)
  );
  Odrv4 odrv_17_17_66246_66142 (
    .I(net_66246),
    .O(net_66142)
  );
  Odrv4 odrv_17_17_66246_66379 (
    .I(net_66246),
    .O(net_66379)
  );
  Odrv4 odrv_17_18_66368_58847 (
    .I(net_66368),
    .O(net_58847)
  );
  Odrv4 odrv_17_18_66368_66391 (
    .I(net_66368),
    .O(net_66391)
  );
  Odrv4 odrv_17_2_64358_68360 (
    .I(net_64358),
    .O(net_68360)
  );
  Odrv4 odrv_17_2_64365_64534 (
    .I(net_64365),
    .O(net_64534)
  );
  Odrv4 odrv_17_3_64519_56992 (
    .I(net_64519),
    .O(net_56992)
  );
  Odrv4 odrv_17_4_64642_68248 (
    .I(net_64642),
    .O(net_68248)
  );
  Odrv4 odrv_17_6_64893_65026 (
    .I(net_64893),
    .O(net_65026)
  );
  Odrv4 odrv_17_7_65016_57486 (
    .I(net_65016),
    .O(net_57486)
  );
  Odrv4 odrv_17_7_65016_64912 (
    .I(net_65016),
    .O(net_64912)
  );
  Odrv4 odrv_17_8_65133_61438 (
    .I(net_65133),
    .O(net_61438)
  );
  Odrv4 odrv_17_8_65134_57607 (
    .I(net_65134),
    .O(net_57607)
  );
  Odrv4 odrv_17_8_65138_57617 (
    .I(net_65138),
    .O(net_57617)
  );
  Odrv4 odrv_17_9_65259_65042 (
    .I(net_65259),
    .O(net_65042)
  );
  Odrv4 odrv_18_0_68185_60431 (
    .I(net_68185),
    .O(net_60431)
  );
  Odrv4 odrv_18_10_69211_72950 (
    .I(net_69211),
    .O(net_72950)
  );
  Odrv4 odrv_18_10_69214_65517 (
    .I(net_69214),
    .O(net_65517)
  );
  Odrv4 odrv_18_10_69216_65521 (
    .I(net_69216),
    .O(net_65521)
  );
  Odrv4 odrv_18_11_69336_61812 (
    .I(net_69336),
    .O(net_61812)
  );
  Odrv4 odrv_18_11_69336_65636 (
    .I(net_69336),
    .O(net_65636)
  );
  Odrv4 odrv_18_11_69336_69357 (
    .I(net_69336),
    .O(net_69357)
  );
  Odrv4 odrv_18_11_69336_73308 (
    .I(net_69336),
    .O(net_73308)
  );
  Odrv4 odrv_18_12_69462_69358 (
    .I(net_69462),
    .O(net_69358)
  );
  Odrv4 odrv_18_13_69579_65884 (
    .I(net_69579),
    .O(net_65884)
  );
  Odrv4 odrv_18_13_69580_62052 (
    .I(net_69580),
    .O(net_62052)
  );
  Odrv4 odrv_18_13_69582_62058 (
    .I(net_69582),
    .O(net_62058)
  );
  Odrv4 odrv_18_13_69583_69367 (
    .I(net_69583),
    .O(net_69367)
  );
  Odrv4 odrv_18_13_69584_62062 (
    .I(net_69584),
    .O(net_62062)
  );
  Odrv4 odrv_18_14_69701_66015 (
    .I(net_69701),
    .O(net_66015)
  );
  Odrv4 odrv_18_14_69703_62175 (
    .I(net_69703),
    .O(net_62175)
  );
  Odrv4 odrv_18_14_69704_62179 (
    .I(net_69704),
    .O(net_62179)
  );
  Odrv4 odrv_18_14_69705_62181 (
    .I(net_69705),
    .O(net_62181)
  );
  Odrv4 odrv_18_14_69706_73320 (
    .I(net_69706),
    .O(net_73320)
  );
  Odrv4 odrv_18_14_69707_69602 (
    .I(net_69707),
    .O(net_69602)
  );
  Odrv4 odrv_18_14_69708_66013 (
    .I(net_69708),
    .O(net_66013)
  );
  Odrv4 odrv_18_16_69948_66253 (
    .I(net_69948),
    .O(net_66253)
  );
  Odrv4 odrv_18_16_69948_69728 (
    .I(net_69948),
    .O(net_69728)
  );
  Odrv4 odrv_18_16_69949_69730 (
    .I(net_69949),
    .O(net_69730)
  );
  Odrv4 odrv_18_16_69952_69736 (
    .I(net_69952),
    .O(net_69736)
  );
  Odrv4 odrv_18_16_69954_69978 (
    .I(net_69954),
    .O(net_69978)
  );
  Odrv4 odrv_18_2_68193_60705 (
    .I(net_68193),
    .O(net_60705)
  );
  Odrv4 odrv_18_2_68193_64529 (
    .I(net_68193),
    .O(net_64529)
  );
  Odrv4 odrv_18_3_68354_68503 (
    .I(net_68354),
    .O(net_68503)
  );
  Odrv4 odrv_18_4_68472_72441 (
    .I(net_68472),
    .O(net_72441)
  );
  Odrv4 odrv_18_4_68473_68618 (
    .I(net_68473),
    .O(net_68618)
  );
  Odrv4 odrv_18_4_68474_68620 (
    .I(net_68474),
    .O(net_68620)
  );
  Odrv4 odrv_18_4_68475_68622 (
    .I(net_68475),
    .O(net_68622)
  );
  Odrv4 odrv_18_4_68476_68624 (
    .I(net_68476),
    .O(net_68624)
  );
  Odrv4 odrv_18_4_68477_72458 (
    .I(net_68477),
    .O(net_72458)
  );
  Odrv4 odrv_18_4_68478_72460 (
    .I(net_68478),
    .O(net_72460)
  );
  Odrv4 odrv_18_5_68594_72560 (
    .I(net_68594),
    .O(net_72560)
  );
  Odrv4 odrv_18_5_68595_72564 (
    .I(net_68595),
    .O(net_72564)
  );
  Odrv4 odrv_18_6_68717_68496 (
    .I(net_68717),
    .O(net_68496)
  );
  Odrv4 odrv_18_6_68721_68504 (
    .I(net_68721),
    .O(net_68504)
  );
  Odrv4 odrv_18_6_68724_72452 (
    .I(net_68724),
    .O(net_72452)
  );
  Odrv4 odrv_18_7_68841_68875 (
    .I(net_68841),
    .O(net_68875)
  );
  Odrv12 odrv_18_7_68841_72435 (
    .I(net_68841),
    .O(net_72435)
  );
  Odrv4 odrv_18_7_68841_72810 (
    .I(net_68841),
    .O(net_72810)
  );
  Odrv4 odrv_18_7_68842_68986 (
    .I(net_68842),
    .O(net_68986)
  );
  Odrv4 odrv_18_7_68842_68987 (
    .I(net_68842),
    .O(net_68987)
  );
  Odrv12 odrv_18_7_68843_45988 (
    .I(net_68843),
    .O(net_45988)
  );
  Odrv4 odrv_18_7_68843_68989 (
    .I(net_68843),
    .O(net_68989)
  );
  Odrv12 odrv_18_7_68844_42156 (
    .I(net_68844),
    .O(net_42156)
  );
  Odrv4 odrv_18_7_68844_61320 (
    .I(net_68844),
    .O(net_61320)
  );
  Odrv4 odrv_18_7_68844_68865 (
    .I(net_68844),
    .O(net_68865)
  );
  Odrv12 odrv_18_7_68845_38326 (
    .I(net_68845),
    .O(net_38326)
  );
  Odrv4 odrv_18_7_68845_61322 (
    .I(net_68845),
    .O(net_61322)
  );
  Odrv4 odrv_18_7_68845_68993 (
    .I(net_68845),
    .O(net_68993)
  );
  Odrv4 odrv_18_7_68846_65150 (
    .I(net_68846),
    .O(net_65150)
  );
  Odrv4 odrv_18_7_68846_68869 (
    .I(net_68846),
    .O(net_68869)
  );
  Odrv4 odrv_18_7_68846_68995 (
    .I(net_68846),
    .O(net_68995)
  );
  Odrv4 odrv_18_7_68847_68743 (
    .I(net_68847),
    .O(net_68743)
  );
  Odrv4 odrv_18_7_68847_68980 (
    .I(net_68847),
    .O(net_68980)
  );
  Odrv4 odrv_18_8_68963_65277 (
    .I(net_68963),
    .O(net_65277)
  );
  Odrv4 odrv_18_8_68963_68996 (
    .I(net_68963),
    .O(net_68996)
  );
  Odrv4 odrv_18_8_68963_72929 (
    .I(net_68963),
    .O(net_72929)
  );
  Odrv4 odrv_18_8_68964_69107 (
    .I(net_68964),
    .O(net_69107)
  );
  Odrv4 odrv_18_8_68964_72702 (
    .I(net_68964),
    .O(net_72702)
  );
  Odrv4 odrv_18_8_68964_72933 (
    .I(net_68964),
    .O(net_72933)
  );
  Odrv4 odrv_18_8_68967_61443 (
    .I(net_68967),
    .O(net_61443)
  );
  Odrv4 odrv_18_8_68968_68752 (
    .I(net_68968),
    .O(net_68752)
  );
  Odrv4 odrv_18_8_68970_61439 (
    .I(net_68970),
    .O(net_61439)
  );
  Odrv4 odrv_18_9_69087_65392 (
    .I(net_69087),
    .O(net_65392)
  );
  Odrv4 odrv_18_9_69089_72829 (
    .I(net_69089),
    .O(net_72829)
  );
  Odrv4 odrv_19_0_72016_64262 (
    .I(net_72016),
    .O(net_64262)
  );
  Odrv4 odrv_19_0_72018_72048 (
    .I(net_72018),
    .O(net_72048)
  );
  Odrv4 odrv_1_10_1967_7771 (
    .I(net_1967),
    .O(net_7771)
  );
  Odrv4 odrv_1_10_1967_8202 (
    .I(net_1967),
    .O(net_8202)
  );
  Odrv4 odrv_1_10_1971_2239 (
    .I(net_1971),
    .O(net_2239)
  );
  Odrv4 odrv_1_10_1971_7915 (
    .I(net_1971),
    .O(net_7915)
  );
  Odrv4 odrv_1_10_1971_8065 (
    .I(net_1971),
    .O(net_8065)
  );
  Odrv4 odrv_1_11_2193_1856 (
    .I(net_2193),
    .O(net_1856)
  );
  Odrv4 odrv_1_11_2193_7920 (
    .I(net_2193),
    .O(net_7920)
  );
  Odrv4 odrv_1_11_2193_8072 (
    .I(net_2193),
    .O(net_8072)
  );
  Odrv4 odrv_1_11_2193_8351 (
    .I(net_2193),
    .O(net_8351)
  );
  Odrv4 odrv_1_11_2196_2291 (
    .I(net_2196),
    .O(net_2291)
  );
  Odrv4 odrv_1_12_2396_8363 (
    .I(net_2396),
    .O(net_8363)
  );
  Odrv4 odrv_1_12_2398_2670 (
    .I(net_2398),
    .O(net_2670)
  );
  Odrv4 odrv_1_12_2400_2657 (
    .I(net_2400),
    .O(net_2657)
  );
  Odrv4 odrv_1_12_2403_8361 (
    .I(net_2403),
    .O(net_8361)
  );
  Odrv4 odrv_1_13_2604_8637 (
    .I(net_2604),
    .O(net_8637)
  );
  Odrv4 odrv_1_13_2605_8641 (
    .I(net_2605),
    .O(net_8641)
  );
  Odrv4 odrv_1_13_2606_8643 (
    .I(net_2606),
    .O(net_8643)
  );
  Odrv4 odrv_1_13_2607_2864 (
    .I(net_2607),
    .O(net_2864)
  );
  Odrv4 odrv_1_13_2608_8647 (
    .I(net_2608),
    .O(net_8647)
  );
  Odrv4 odrv_1_13_2609_2868 (
    .I(net_2609),
    .O(net_2868)
  );
  Odrv4 odrv_1_13_2610_2870 (
    .I(net_2610),
    .O(net_2870)
  );
  Odrv4 odrv_1_13_2611_2872 (
    .I(net_2611),
    .O(net_2872)
  );
  Odrv4 odrv_1_14_2813_2493 (
    .I(net_2813),
    .O(net_2493)
  );
  Odrv4 odrv_1_14_2815_2497 (
    .I(net_2815),
    .O(net_2497)
  );
  Odrv4 odrv_1_14_2818_2503 (
    .I(net_2818),
    .O(net_2503)
  );
  Odrv4 odrv_1_14_2820_8505 (
    .I(net_2820),
    .O(net_8505)
  );
  Odrv4 odrv_1_16_3251_9082 (
    .I(net_3251),
    .O(net_9082)
  );
  Odrv4 odrv_1_17_3459_8802 (
    .I(net_3459),
    .O(net_8802)
  );
  Odrv4 odrv_1_17_3463_3348 (
    .I(net_3463),
    .O(net_3348)
  );
  Odrv4 odrv_1_1_107_6871 (
    .I(net_107),
    .O(net_6871)
  );
  Odrv4 odrv_1_1_107_6889 (
    .I(net_107),
    .O(net_6889)
  );
  Odrv4 odrv_1_1_108_292 (
    .I(net_108),
    .O(net_292)
  );
  Odrv4 odrv_1_21_4315_3976 (
    .I(net_4315),
    .O(net_3976)
  );
  Odrv4 odrv_1_22_4545_4423 (
    .I(net_4545),
    .O(net_4423)
  );
  Odrv4 odrv_1_2_122_523 (
    .I(net_122),
    .O(net_523)
  );
  Odrv4 odrv_1_3_453_788 (
    .I(net_453),
    .O(net_788)
  );
  Odrv4 odrv_1_3_454_761 (
    .I(net_454),
    .O(net_761)
  );
  Odrv4 odrv_1_3_455_7177 (
    .I(net_455),
    .O(net_7177)
  );
  Odrv4 odrv_1_3_456_7169 (
    .I(net_456),
    .O(net_7169)
  );
  Odrv4 odrv_1_5_905_7032 (
    .I(net_905),
    .O(net_7032)
  );
  Odrv4 odrv_1_5_906_1027 (
    .I(net_906),
    .O(net_1027)
  );
  Odrv4 odrv_1_5_906_1223 (
    .I(net_906),
    .O(net_1223)
  );
  Odrv4 odrv_1_5_907_1225 (
    .I(net_907),
    .O(net_1225)
  );
  Odrv4 odrv_1_5_908_1181 (
    .I(net_908),
    .O(net_1181)
  );
  Odrv4 odrv_1_5_909_1017 (
    .I(net_909),
    .O(net_1017)
  );
  Odrv4 odrv_1_5_909_571 (
    .I(net_909),
    .O(net_571)
  );
  Odrv4 odrv_1_5_912_1201 (
    .I(net_912),
    .O(net_1201)
  );
  Odrv4 odrv_1_5_912_1236 (
    .I(net_912),
    .O(net_1236)
  );
  Odrv12 odrv_1_6_1133_7459 (
    .I(net_1133),
    .O(net_7459)
  );
  Odrv4 odrv_1_6_1134_1436 (
    .I(net_1134),
    .O(net_1436)
  );
  Odrv4 odrv_1_6_1136_1440 (
    .I(net_1136),
    .O(net_1440)
  );
  Odrv4 odrv_1_8_1547_1851 (
    .I(net_1547),
    .O(net_1851)
  );
  Odrv4 odrv_1_8_1548_1853 (
    .I(net_1548),
    .O(net_1853)
  );
  Odrv4 odrv_1_8_1549_7904 (
    .I(net_1549),
    .O(net_7904)
  );
  Odrv4 odrv_1_8_1551_1647 (
    .I(net_1551),
    .O(net_1647)
  );
  Odrv4 odrv_1_9_1753_1858 (
    .I(net_1753),
    .O(net_1858)
  );
  Odrv4 odrv_1_9_1753_2071 (
    .I(net_1753),
    .O(net_2071)
  );
  Odrv4 odrv_1_9_1754_1860 (
    .I(net_1754),
    .O(net_1860)
  );
  Odrv4 odrv_1_9_1755_2076 (
    .I(net_1755),
    .O(net_2076)
  );
  Odrv4 odrv_1_9_1756_2078 (
    .I(net_1756),
    .O(net_2078)
  );
  Odrv4 odrv_1_9_1757_1850 (
    .I(net_1757),
    .O(net_1850)
  );
  Odrv4 odrv_1_9_1757_8066 (
    .I(net_1757),
    .O(net_8066)
  );
  Odrv4 odrv_1_9_1759_7918 (
    .I(net_1759),
    .O(net_7918)
  );
  Odrv4 odrv_1_9_1759_8070 (
    .I(net_1759),
    .O(net_8070)
  );
  Odrv4 odrv_20_10_76655_73175 (
    .I(net_76655),
    .O(net_73175)
  );
  Odrv4 odrv_20_10_76656_73179 (
    .I(net_76656),
    .O(net_73179)
  );
  Odrv4 odrv_20_11_76760_73306 (
    .I(net_76760),
    .O(net_73306)
  );
  Odrv4 odrv_20_12_76857_76710 (
    .I(net_76857),
    .O(net_76710)
  );
  Odrv4 odrv_20_14_77062_69841 (
    .I(net_77062),
    .O(net_69841)
  );
  Odrv4 odrv_20_2_75801_68361 (
    .I(net_75801),
    .O(net_68361)
  );
  Odrv4 odrv_20_2_75806_68363 (
    .I(net_75806),
    .O(net_68363)
  );
  Odrv4 odrv_20_3_75940_68488 (
    .I(net_75940),
    .O(net_68488)
  );
  Odrv4 odrv_20_3_75942_68492 (
    .I(net_75942),
    .O(net_68492)
  );
  Odrv4 odrv_20_3_75943_72320 (
    .I(net_75943),
    .O(net_72320)
  );
  Odrv4 odrv_20_3_75944_68486 (
    .I(net_75944),
    .O(net_68486)
  );
  Odrv4 odrv_20_4_76040_76192 (
    .I(net_76040),
    .O(net_76192)
  );
  Odrv4 odrv_20_4_76040_79241 (
    .I(net_76040),
    .O(net_79241)
  );
  Odrv4 odrv_20_5_76141_76292 (
    .I(net_76141),
    .O(net_76292)
  );
  Odrv4 odrv_20_5_76142_79595 (
    .I(net_76142),
    .O(net_79595)
  );
  Odrv4 odrv_20_5_76143_68730 (
    .I(net_76143),
    .O(net_68730)
  );
  Odrv4 odrv_20_5_76144_68734 (
    .I(net_76144),
    .O(net_68734)
  );
  Odrv4 odrv_20_5_76145_68736 (
    .I(net_76145),
    .O(net_68736)
  );
  Odrv4 odrv_20_5_76146_68738 (
    .I(net_76146),
    .O(net_68738)
  );
  Odrv4 odrv_20_5_76147_72566 (
    .I(net_76147),
    .O(net_72566)
  );
  Odrv4 odrv_20_5_76148_68732 (
    .I(net_76148),
    .O(net_68732)
  );
  Odrv4 odrv_20_6_76243_72693 (
    .I(net_76243),
    .O(net_72693)
  );
  Odrv4 odrv_20_6_76247_68859 (
    .I(net_76247),
    .O(net_68859)
  );
  Odrv4 odrv_20_6_76248_76300 (
    .I(net_76248),
    .O(net_76300)
  );
  Odrv4 odrv_20_7_76350_68984 (
    .I(net_76350),
    .O(net_68984)
  );
  Odrv4 odrv_20_8_76453_76506 (
    .I(net_76453),
    .O(net_76506)
  );
  Odrv4 odrv_20_8_76453_76592 (
    .I(net_76453),
    .O(net_76592)
  );
  Odrv4 odrv_20_9_76552_76511 (
    .I(net_76552),
    .O(net_76511)
  );
  Odrv4 odrv_20_9_76553_80093 (
    .I(net_76553),
    .O(net_80093)
  );
  Odrv4 odrv_20_9_76554_69230 (
    .I(net_76554),
    .O(net_69230)
  );
  Odrv4 odrv_21_10_80071_84037 (
    .I(net_80071),
    .O(net_84037)
  );
  Odrv4 odrv_21_10_80072_84041 (
    .I(net_80072),
    .O(net_84041)
  );
  Odrv4 odrv_21_10_80075_73182 (
    .I(net_80075),
    .O(net_73182)
  );
  Odrv4 odrv_21_3_79210_83176 (
    .I(net_79210),
    .O(net_83176)
  );
  Odrv4 odrv_21_3_79212_72315 (
    .I(net_79212),
    .O(net_72315)
  );
  Odrv4 odrv_21_3_79217_72317 (
    .I(net_79217),
    .O(net_72317)
  );
  Odrv4 odrv_21_4_79333_79475 (
    .I(net_79333),
    .O(net_79475)
  );
  Odrv4 odrv_21_4_79334_79477 (
    .I(net_79334),
    .O(net_79477)
  );
  Odrv4 odrv_21_4_79335_72438 (
    .I(net_79335),
    .O(net_72438)
  );
  Odrv4 odrv_21_4_79338_72446 (
    .I(net_79338),
    .O(net_72446)
  );
  Odrv4 odrv_21_4_79340_72440 (
    .I(net_79340),
    .O(net_72440)
  );
  Odrv4 odrv_21_5_79458_72561 (
    .I(net_79458),
    .O(net_72561)
  );
  Odrv4 odrv_21_5_79460_72567 (
    .I(net_79460),
    .O(net_72567)
  );
  Odrv4 odrv_21_5_79462_72571 (
    .I(net_79462),
    .O(net_72571)
  );
  Odrv4 odrv_21_6_79583_72690 (
    .I(net_79583),
    .O(net_72690)
  );
  Odrv4 odrv_21_6_79584_72692 (
    .I(net_79584),
    .O(net_72692)
  );
  Odrv4 odrv_21_6_79586_79719 (
    .I(net_79586),
    .O(net_79719)
  );
  Odrv4 odrv_21_7_79705_72811 (
    .I(net_79705),
    .O(net_72811)
  );
  Odrv4 odrv_21_7_79709_72809 (
    .I(net_79709),
    .O(net_72809)
  );
  Odrv12 odrv_21_8_79827_61432 (
    .I(net_79827),
    .O(net_61432)
  );
  Odrv12 odrv_21_8_79828_57603 (
    .I(net_79828),
    .O(net_57603)
  );
  Odrv4 odrv_21_8_79829_72936 (
    .I(net_79829),
    .O(net_72936)
  );
  Odrv4 odrv_21_8_79830_79852 (
    .I(net_79830),
    .O(net_79852)
  );
  Odrv4 odrv_21_8_79831_72940 (
    .I(net_79831),
    .O(net_72940)
  );
  Odrv4 odrv_21_9_79949_79855 (
    .I(net_79949),
    .O(net_79855)
  );
  Odrv4 odrv_21_9_79950_80094 (
    .I(net_79950),
    .O(net_80094)
  );
  Odrv4 odrv_22_10_83902_80216 (
    .I(net_83902),
    .O(net_80216)
  );
  Odrv4 odrv_22_10_83902_83681 (
    .I(net_83902),
    .O(net_83681)
  );
  Odrv4 odrv_22_10_83902_83935 (
    .I(net_83902),
    .O(net_83935)
  );
  Odrv12 odrv_22_10_83902_87375 (
    .I(net_83902),
    .O(net_87375)
  );
  Odrv4 odrv_22_10_83902_87639 (
    .I(net_83902),
    .O(net_87639)
  );
  Odrv4 odrv_22_10_83902_87765 (
    .I(net_83902),
    .O(net_87765)
  );
  Odrv4 odrv_22_3_83045_87017 (
    .I(net_83045),
    .O(net_87017)
  );
  Odrv12 odrv_22_4_83166_64771 (
    .I(net_83166),
    .O(net_64771)
  );
  Odrv4 odrv_22_5_83287_79601 (
    .I(net_83287),
    .O(net_79601)
  );
  Odrv4 odrv_22_5_83290_76290 (
    .I(net_83290),
    .O(net_76290)
  );
  Odrv4 odrv_22_5_83294_83427 (
    .I(net_83294),
    .O(net_83427)
  );
  Odrv4 odrv_22_6_83416_83546 (
    .I(net_83416),
    .O(net_83546)
  );
  Odrv4 odrv_23_0_86709_86737 (
    .I(net_86709),
    .O(net_86737)
  );
  Odrv4 odrv_23_0_86709_86745 (
    .I(net_86709),
    .O(net_86745)
  );
  Odrv4 odrv_23_5_87122_79598 (
    .I(net_87122),
    .O(net_79598)
  );
  Odrv4 odrv_23_5_87123_87145 (
    .I(net_87123),
    .O(net_87145)
  );
  Odrv4 odrv_23_8_87494_83799 (
    .I(net_87494),
    .O(net_83799)
  );
  Odrv4 odrv_23_9_87613_80088 (
    .I(net_87613),
    .O(net_80088)
  );
  Odrv4 odrv_25_10_100050_95258 (
    .I(net_100050),
    .O(net_95258)
  );
  Odrv4 odrv_25_10_100051_91701 (
    .I(net_100051),
    .O(net_91701)
  );
  Odrv4 odrv_25_10_100052_87869 (
    .I(net_100052),
    .O(net_87869)
  );
  Odrv4 odrv_25_10_100053_87873 (
    .I(net_100053),
    .O(net_87873)
  );
  Odrv4 odrv_25_10_100054_91699 (
    .I(net_100054),
    .O(net_91699)
  );
  Odrv4 odrv_25_10_100055_91703 (
    .I(net_100055),
    .O(net_91703)
  );
  Odrv4 odrv_25_10_100056_91705 (
    .I(net_100056),
    .O(net_91705)
  );
  Odrv4 odrv_25_10_100057_87871 (
    .I(net_100057),
    .O(net_87871)
  );
  Odrv4 odrv_25_11_100200_87992 (
    .I(net_100200),
    .O(net_87992)
  );
  Odrv4 odrv_25_11_100201_95545 (
    .I(net_100201),
    .O(net_95545)
  );
  Odrv4 odrv_25_11_100202_95405 (
    .I(net_100202),
    .O(net_95405)
  );
  Odrv4 odrv_25_11_100203_95407 (
    .I(net_100203),
    .O(net_95407)
  );
  Odrv4 odrv_25_11_100204_95535 (
    .I(net_100204),
    .O(net_95535)
  );
  Odrv4 odrv_25_11_100205_87994 (
    .I(net_100205),
    .O(net_87994)
  );
  Odrv4 odrv_25_11_100206_95397 (
    .I(net_100206),
    .O(net_95397)
  );
  Odrv4 odrv_25_11_100207_100240 (
    .I(net_100207),
    .O(net_100240)
  );
  Odrv4 odrv_25_12_100352_95678 (
    .I(net_100352),
    .O(net_95678)
  );
  Odrv4 odrv_25_12_100353_95538 (
    .I(net_100353),
    .O(net_95538)
  );
  Odrv4 odrv_25_12_100354_95682 (
    .I(net_100354),
    .O(net_95682)
  );
  Odrv4 odrv_25_12_100355_95542 (
    .I(net_100355),
    .O(net_95542)
  );
  Odrv4 odrv_25_12_100356_88121 (
    .I(net_100356),
    .O(net_88121)
  );
  Odrv4 odrv_25_12_100357_95546 (
    .I(net_100357),
    .O(net_95546)
  );
  Odrv4 odrv_25_12_100358_91951 (
    .I(net_100358),
    .O(net_91951)
  );
  Odrv4 odrv_25_12_100359_88117 (
    .I(net_100359),
    .O(net_88117)
  );
  Odrv4 odrv_25_13_100504_95675 (
    .I(net_100504),
    .O(net_95675)
  );
  Odrv4 odrv_25_13_100505_95677 (
    .I(net_100505),
    .O(net_95677)
  );
  Odrv4 odrv_25_13_100506_96090 (
    .I(net_100506),
    .O(net_96090)
  );
  Odrv4 odrv_25_13_100507_88242 (
    .I(net_100507),
    .O(net_88242)
  );
  Odrv4 odrv_25_13_100508_88244 (
    .I(net_100508),
    .O(net_88244)
  );
  Odrv4 odrv_25_13_100509_95685 (
    .I(net_100509),
    .O(net_95685)
  );
  Odrv4 odrv_25_13_100510_88248 (
    .I(net_100510),
    .O(net_88248)
  );
  Odrv4 odrv_25_13_100511_92076 (
    .I(net_100511),
    .O(net_92076)
  );
  Odrv4 odrv_25_5_99270_91094 (
    .I(net_99270),
    .O(net_91094)
  );
  Odrv4 odrv_25_5_99271_94851 (
    .I(net_99271),
    .O(net_94851)
  );
  Odrv4 odrv_25_5_99272_87254 (
    .I(net_99272),
    .O(net_87254)
  );
  Odrv4 odrv_25_5_99273_87258 (
    .I(net_99273),
    .O(net_87258)
  );
  Odrv4 odrv_25_5_99274_91084 (
    .I(net_99274),
    .O(net_91084)
  );
  Odrv4 odrv_25_5_99275_87262 (
    .I(net_99275),
    .O(net_87262)
  );
  Odrv4 odrv_25_5_99276_87264 (
    .I(net_99276),
    .O(net_87264)
  );
  Odrv4 odrv_25_5_99277_87256 (
    .I(net_99277),
    .O(net_87256)
  );
  Odrv4 odrv_25_6_99420_87377 (
    .I(net_99420),
    .O(net_87377)
  );
  Odrv4 odrv_25_6_99421_95109 (
    .I(net_99421),
    .O(net_95109)
  );
  Odrv4 odrv_25_6_99422_87383 (
    .I(net_99422),
    .O(net_87383)
  );
  Odrv4 odrv_25_6_99423_99458 (
    .I(net_99423),
    .O(net_99458)
  );
  Odrv4 odrv_25_6_99424_95107 (
    .I(net_99424),
    .O(net_95107)
  );
  Odrv4 odrv_25_6_99425_94986 (
    .I(net_99425),
    .O(net_94986)
  );
  Odrv4 odrv_25_6_99426_91217 (
    .I(net_99426),
    .O(net_91217)
  );
  Odrv4 odrv_25_6_99427_91209 (
    .I(net_99427),
    .O(net_91209)
  );
  Odrv4 odrv_25_7_99572_94841 (
    .I(net_99572),
    .O(net_94841)
  );
  Odrv4 odrv_25_7_99573_94843 (
    .I(net_99573),
    .O(net_94843)
  );
  Odrv4 odrv_25_7_99574_94987 (
    .I(net_99574),
    .O(net_94987)
  );
  Odrv4 odrv_25_7_99575_95259 (
    .I(net_99575),
    .O(net_95259)
  );
  Odrv4 odrv_25_7_99576_91330 (
    .I(net_99576),
    .O(net_91330)
  );
  Odrv4 odrv_25_7_99577_87508 (
    .I(net_99577),
    .O(net_87508)
  );
  Odrv4 odrv_25_7_99578_87510 (
    .I(net_99578),
    .O(net_87510)
  );
  Odrv4 odrv_25_7_99579_87502 (
    .I(net_99579),
    .O(net_87502)
  );
  Odrv4 odrv_25_8_99724_91463 (
    .I(net_99724),
    .O(net_91463)
  );
  Odrv4 odrv_25_8_99725_95124 (
    .I(net_99725),
    .O(net_95124)
  );
  Odrv4 odrv_25_8_99726_94984 (
    .I(net_99726),
    .O(net_94984)
  );
  Odrv4 odrv_25_8_99727_95128 (
    .I(net_99727),
    .O(net_95128)
  );
  Odrv4 odrv_25_8_99728_87629 (
    .I(net_99728),
    .O(net_87629)
  );
  Odrv4 odrv_25_8_99729_87631 (
    .I(net_99729),
    .O(net_87631)
  );
  Odrv4 odrv_25_8_99730_87633 (
    .I(net_99730),
    .O(net_87633)
  );
  Odrv4 odrv_25_8_99731_95264 (
    .I(net_99731),
    .O(net_95264)
  );
  Odrv4 odrv_2_10_8039_12525 (
    .I(net_8039),
    .O(net_12525)
  );
  Odrv4 odrv_2_10_8042_2248 (
    .I(net_8042),
    .O(net_2248)
  );
  Odrv4 odrv_2_11_8188_7923 (
    .I(net_8188),
    .O(net_7923)
  );
  Odrv4 odrv_2_11_8191_12530 (
    .I(net_8191),
    .O(net_12530)
  );
  Odrv4 odrv_2_11_8191_12658 (
    .I(net_8191),
    .O(net_12658)
  );
  Odrv4 odrv_2_12_8338_12653 (
    .I(net_8338),
    .O(net_12653)
  );
  Odrv4 odrv_2_13_8480_12887 (
    .I(net_8480),
    .O(net_12887)
  );
  Odrv4 odrv_2_13_8481_12889 (
    .I(net_8481),
    .O(net_12889)
  );
  Odrv4 odrv_2_13_8483_12534 (
    .I(net_8483),
    .O(net_12534)
  );
  Odrv4 odrv_2_13_8483_12883 (
    .I(net_8483),
    .O(net_12883)
  );
  Odrv4 odrv_2_13_8483_2873 (
    .I(net_8483),
    .O(net_2873)
  );
  Odrv4 odrv_2_13_8483_8219 (
    .I(net_8483),
    .O(net_8219)
  );
  Odrv4 odrv_2_13_8484_8355 (
    .I(net_8484),
    .O(net_8355)
  );
  Odrv4 odrv_2_14_8626_12903 (
    .I(net_8626),
    .O(net_12903)
  );
  Odrv4 odrv_2_14_8627_3092 (
    .I(net_8627),
    .O(net_3092)
  );
  Odrv4 odrv_2_14_8628_8362 (
    .I(net_8628),
    .O(net_8362)
  );
  Odrv4 odrv_2_14_8629_8364 (
    .I(net_8629),
    .O(net_8364)
  );
  Odrv4 odrv_2_14_8630_13006 (
    .I(net_8630),
    .O(net_13006)
  );
  Odrv4 odrv_2_14_8631_8785 (
    .I(net_8631),
    .O(net_8785)
  );
  Odrv4 odrv_2_14_8632_12899 (
    .I(net_8632),
    .O(net_12899)
  );
  Odrv4 odrv_2_15_8777_13129 (
    .I(net_8777),
    .O(net_13129)
  );
  Odrv4 odrv_2_15_8779_8936 (
    .I(net_8779),
    .O(net_8936)
  );
  Odrv4 odrv_2_19_9363_9097 (
    .I(net_9363),
    .O(net_9097)
  );
  Odrv4 odrv_2_1_6678_6886 (
    .I(net_6678),
    .O(net_6886)
  );
  Odrv4 odrv_2_21_9655_9387 (
    .I(net_9655),
    .O(net_9387)
  );
  Odrv4 odrv_2_2_6825_11528 (
    .I(net_6825),
    .O(net_11528)
  );
  Odrv4 odrv_2_2_6828_11536 (
    .I(net_6828),
    .O(net_11536)
  );
  Odrv4 odrv_2_2_6828_11543 (
    .I(net_6828),
    .O(net_11543)
  );
  Odrv4 odrv_2_2_6828_7023 (
    .I(net_6828),
    .O(net_7023)
  );
  Odrv4 odrv_2_2_6829_11538 (
    .I(net_6829),
    .O(net_11538)
  );
  Odrv4 odrv_2_2_6829_7036 (
    .I(net_6829),
    .O(net_7036)
  );
  Odrv4 odrv_2_3_7010_11421 (
    .I(net_7010),
    .O(net_11421)
  );
  Odrv4 odrv_2_3_7011_11423 (
    .I(net_7011),
    .O(net_11423)
  );
  Odrv4 odrv_2_4_7160_11776 (
    .I(net_7160),
    .O(net_11776)
  );
  Odrv4 odrv_2_4_7160_6891 (
    .I(net_7160),
    .O(net_6891)
  );
  Odrv4 odrv_2_5_7302_1224 (
    .I(net_7302),
    .O(net_1224)
  );
  Odrv4 odrv_2_5_7302_7335 (
    .I(net_7302),
    .O(net_7335)
  );
  Odrv4 odrv_2_5_7305_11912 (
    .I(net_7305),
    .O(net_11912)
  );
  Odrv4 odrv_2_5_7308_11790 (
    .I(net_7308),
    .O(net_11790)
  );
  Odrv4 odrv_2_5_7308_7179 (
    .I(net_7308),
    .O(net_7179)
  );
  Odrv4 odrv_2_6_7450_1386 (
    .I(net_7450),
    .O(net_1386)
  );
  Odrv4 odrv_2_6_7451_11795 (
    .I(net_7451),
    .O(net_11795)
  );
  Odrv4 odrv_2_6_7451_7619 (
    .I(net_7451),
    .O(net_7619)
  );
  Odrv4 odrv_2_6_7454_12022 (
    .I(net_7454),
    .O(net_12022)
  );
  Odrv4 odrv_2_6_7455_11787 (
    .I(net_7455),
    .O(net_11787)
  );
  Odrv4 odrv_2_7_7597_11788 (
    .I(net_7597),
    .O(net_11788)
  );
  Odrv4 odrv_2_8_7743_12163 (
    .I(net_7743),
    .O(net_12163)
  );
  Odrv4 odrv_2_8_7744_12165 (
    .I(net_7744),
    .O(net_12165)
  );
  Odrv4 odrv_2_8_7746_12274 (
    .I(net_7746),
    .O(net_12274)
  );
  Odrv4 odrv_2_8_7747_12276 (
    .I(net_7747),
    .O(net_12276)
  );
  Odrv4 odrv_2_9_7893_12166 (
    .I(net_7893),
    .O(net_12166)
  );
  Odrv4 odrv_2_9_7893_12404 (
    .I(net_7893),
    .O(net_12404)
  );
  Odrv4 odrv_2_9_7893_8052 (
    .I(net_7893),
    .O(net_8052)
  );
  Odrv4 odrv_2_9_7896_12156 (
    .I(net_7896),
    .O(net_12156)
  );
  Odrv4 odrv_2_9_7896_7767 (
    .I(net_7896),
    .O(net_7767)
  );
  Odrv4 odrv_2_9_7896_8050 (
    .I(net_7896),
    .O(net_8050)
  );
  Odrv4 odrv_2_9_7897_12284 (
    .I(net_7897),
    .O(net_12284)
  );
  Odrv4 odrv_2_9_7897_8071 (
    .I(net_7897),
    .O(net_8071)
  );
  Odrv4 odrv_3_10_12379_12160 (
    .I(net_12379),
    .O(net_12160)
  );
  Odrv4 odrv_3_10_12379_16349 (
    .I(net_12379),
    .O(net_16349)
  );
  Odrv4 odrv_3_10_12383_16236 (
    .I(net_12383),
    .O(net_16236)
  );
  Odrv4 odrv_3_11_12500_16109 (
    .I(net_12500),
    .O(net_16109)
  );
  Odrv4 odrv_3_11_12500_16363 (
    .I(net_12500),
    .O(net_16363)
  );
  Odrv4 odrv_3_11_12501_12407 (
    .I(net_12501),
    .O(net_12407)
  );
  Odrv4 odrv_3_11_12501_16111 (
    .I(net_12501),
    .O(net_16111)
  );
  Odrv4 odrv_3_11_12503_12411 (
    .I(net_12503),
    .O(net_12411)
  );
  Odrv4 odrv_3_11_12503_16115 (
    .I(net_12503),
    .O(net_16115)
  );
  Odrv4 odrv_3_11_12505_16357 (
    .I(net_12505),
    .O(net_16357)
  );
  Odrv4 odrv_3_11_12505_2489 (
    .I(net_12505),
    .O(net_2489)
  );
  Odrv4 odrv_3_11_12506_16359 (
    .I(net_12506),
    .O(net_16359)
  );
  Odrv4 odrv_3_11_12506_2491 (
    .I(net_12506),
    .O(net_2491)
  );
  Odrv4 odrv_3_13_12747_16716 (
    .I(net_12747),
    .O(net_16716)
  );
  Odrv4 odrv_3_13_12748_12892 (
    .I(net_12748),
    .O(net_12892)
  );
  Odrv4 odrv_3_13_12749_12884 (
    .I(net_12749),
    .O(net_12884)
  );
  Odrv4 odrv_3_13_12750_16722 (
    .I(net_12750),
    .O(net_16722)
  );
  Odrv4 odrv_3_13_12751_16714 (
    .I(net_12751),
    .O(net_16714)
  );
  Odrv4 odrv_3_13_12752_12882 (
    .I(net_12752),
    .O(net_12882)
  );
  Odrv4 odrv_3_14_12872_12654 (
    .I(net_12872),
    .O(net_12654)
  );
  Odrv4 odrv_3_14_12873_12894 (
    .I(net_12873),
    .O(net_12894)
  );
  Odrv4 odrv_3_14_12875_12770 (
    .I(net_12875),
    .O(net_12770)
  );
  Odrv4 odrv_3_14_12876_16604 (
    .I(net_12876),
    .O(net_16604)
  );
  Odrv4 odrv_3_15_12993_16731 (
    .I(net_12993),
    .O(net_16731)
  );
  Odrv4 odrv_3_15_12994_12775 (
    .I(net_12994),
    .O(net_12775)
  );
  Odrv4 odrv_3_15_12995_16607 (
    .I(net_12995),
    .O(net_16607)
  );
  Odrv4 odrv_3_15_12996_12779 (
    .I(net_12996),
    .O(net_12779)
  );
  Odrv4 odrv_3_15_12997_12781 (
    .I(net_12997),
    .O(net_12781)
  );
  Odrv4 odrv_3_15_12998_16725 (
    .I(net_12998),
    .O(net_16725)
  );
  Odrv4 odrv_3_15_12999_12895 (
    .I(net_12999),
    .O(net_12895)
  );
  Odrv4 odrv_3_16_13117_12898 (
    .I(net_13117),
    .O(net_12898)
  );
  Odrv4 odrv_3_16_13118_12900 (
    .I(net_13118),
    .O(net_12900)
  );
  Odrv4 odrv_3_16_13121_13016 (
    .I(net_13121),
    .O(net_13016)
  );
  Odrv4 odrv_3_17_13238_13017 (
    .I(net_13238),
    .O(net_13017)
  );
  Odrv4 odrv_3_17_13245_13141 (
    .I(net_13245),
    .O(net_13141)
  );
  Odrv4 odrv_3_18_13361_16970 (
    .I(net_13361),
    .O(net_16970)
  );
  Odrv4 odrv_3_18_13365_13148 (
    .I(net_13365),
    .O(net_13148)
  );
  Odrv4 odrv_3_18_13366_16980 (
    .I(net_13366),
    .O(net_16980)
  );
  Odrv4 odrv_3_18_13367_17094 (
    .I(net_13367),
    .O(net_17094)
  );
  Odrv4 odrv_3_18_13368_13264 (
    .I(net_13368),
    .O(net_13264)
  );
  Odrv4 odrv_3_19_13486_17097 (
    .I(net_13486),
    .O(net_17097)
  );
  Odrv4 odrv_3_1_11230_11378 (
    .I(net_11230),
    .O(net_11378)
  );
  Odrv4 odrv_3_1_11231_11380 (
    .I(net_11231),
    .O(net_11380)
  );
  Odrv4 odrv_3_1_11232_15208 (
    .I(net_11232),
    .O(net_15208)
  );
  Odrv4 odrv_3_1_11235_11370 (
    .I(net_11235),
    .O(net_11370)
  );
  Odrv4 odrv_3_1_11235_15234 (
    .I(net_11235),
    .O(net_15234)
  );
  Odrv4 odrv_3_1_11235_250 (
    .I(net_11235),
    .O(net_250)
  );
  Odrv4 odrv_3_1_11236_11374 (
    .I(net_11236),
    .O(net_11374)
  );
  Odrv4 odrv_3_20_13608_13388 (
    .I(net_13608),
    .O(net_13388)
  );
  Odrv4 odrv_3_21_13735_13519 (
    .I(net_13735),
    .O(net_13519)
  );
  Odrv4 odrv_3_21_13736_13631 (
    .I(net_13736),
    .O(net_13631)
  );
  Odrv4 odrv_3_2_11359_15365 (
    .I(net_11359),
    .O(net_15365)
  );
  Odrv4 odrv_3_2_11361_15369 (
    .I(net_11361),
    .O(net_15369)
  );
  Odrv4 odrv_3_2_11363_15229 (
    .I(net_11363),
    .O(net_15229)
  );
  Odrv4 odrv_3_2_11364_15249 (
    .I(net_11364),
    .O(net_15249)
  );
  Odrv4 odrv_3_3_11518_15488 (
    .I(net_11518),
    .O(net_15488)
  );
  Odrv4 odrv_3_3_11519_15490 (
    .I(net_11519),
    .O(net_15490)
  );
  Odrv4 odrv_3_3_11520_11667 (
    .I(net_11520),
    .O(net_11667)
  );
  Odrv4 odrv_3_4_11639_11672 (
    .I(net_11639),
    .O(net_11672)
  );
  Odrv4 odrv_3_4_11639_15242 (
    .I(net_11639),
    .O(net_15242)
  );
  Odrv4 odrv_3_4_11641_11417 (
    .I(net_11641),
    .O(net_11417)
  );
  Odrv4 odrv_3_4_11641_11548 (
    .I(net_11641),
    .O(net_11548)
  );
  Odrv4 odrv_3_4_11641_15247 (
    .I(net_11641),
    .O(net_15247)
  );
  Odrv4 odrv_3_4_11645_11668 (
    .I(net_11645),
    .O(net_11668)
  );
  Odrv4 odrv_3_4_11645_11775 (
    .I(net_11645),
    .O(net_11775)
  );
  Odrv4 odrv_3_5_11762_11541 (
    .I(net_11762),
    .O(net_11541)
  );
  Odrv4 odrv_3_5_11762_15625 (
    .I(net_11762),
    .O(net_15625)
  );
  Odrv4 odrv_3_5_11762_7471 (
    .I(net_11762),
    .O(net_7471)
  );
  Odrv4 odrv_3_5_11763_7463 (
    .I(net_11763),
    .O(net_7463)
  );
  Odrv4 odrv_3_5_11767_7465 (
    .I(net_11767),
    .O(net_7465)
  );
  Odrv4 odrv_3_5_11769_7469 (
    .I(net_11769),
    .O(net_7469)
  );
  Odrv4 odrv_3_6_11888_11796 (
    .I(net_11888),
    .O(net_11796)
  );
  Odrv4 odrv_3_6_11889_15861 (
    .I(net_11889),
    .O(net_15861)
  );
  Odrv4 odrv_3_6_11891_12021 (
    .I(net_11891),
    .O(net_12021)
  );
  Odrv4 odrv_3_7_12010_11917 (
    .I(net_12010),
    .O(net_11917)
  );
  Odrv4 odrv_3_7_12011_11919 (
    .I(net_12011),
    .O(net_11919)
  );
  Odrv4 odrv_3_7_12013_7759 (
    .I(net_12013),
    .O(net_7759)
  );
  Odrv4 odrv_3_8_12131_12164 (
    .I(net_12131),
    .O(net_12164)
  );
  Odrv4 odrv_3_8_12133_12277 (
    .I(net_12133),
    .O(net_12277)
  );
  Odrv4 odrv_3_8_12138_12288 (
    .I(net_12138),
    .O(net_12288)
  );
  Odrv4 odrv_4_10_16208_16241 (
    .I(net_16208),
    .O(net_16241)
  );
  Odrv4 odrv_4_10_16209_16243 (
    .I(net_16209),
    .O(net_16243)
  );
  Odrv4 odrv_4_10_16210_16354 (
    .I(net_16210),
    .O(net_16354)
  );
  Odrv4 odrv_4_10_16211_16346 (
    .I(net_16211),
    .O(net_16346)
  );
  Odrv4 odrv_4_10_16212_16233 (
    .I(net_16212),
    .O(net_16233)
  );
  Odrv4 odrv_4_10_16213_12516 (
    .I(net_16213),
    .O(net_12516)
  );
  Odrv4 odrv_4_10_16214_16237 (
    .I(net_16214),
    .O(net_16237)
  );
  Odrv4 odrv_4_10_16215_20197 (
    .I(net_16215),
    .O(net_20197)
  );
  Odrv4 odrv_4_11_16331_16364 (
    .I(net_16331),
    .O(net_16364)
  );
  Odrv4 odrv_4_11_16332_16366 (
    .I(net_16332),
    .O(net_16366)
  );
  Odrv4 odrv_4_11_16333_16478 (
    .I(net_16333),
    .O(net_16478)
  );
  Odrv4 odrv_4_11_16334_16116 (
    .I(net_16334),
    .O(net_16116)
  );
  Odrv4 odrv_4_11_16334_16242 (
    .I(net_16334),
    .O(net_16242)
  );
  Odrv4 odrv_4_11_16335_16118 (
    .I(net_16335),
    .O(net_16118)
  );
  Odrv4 odrv_4_11_16335_20186 (
    .I(net_16335),
    .O(net_20186)
  );
  Odrv4 odrv_4_11_16336_20316 (
    .I(net_16336),
    .O(net_20316)
  );
  Odrv4 odrv_4_11_16337_16360 (
    .I(net_16337),
    .O(net_16360)
  );
  Odrv4 odrv_4_11_16337_8354 (
    .I(net_16337),
    .O(net_8354)
  );
  Odrv4 odrv_4_11_16338_16362 (
    .I(net_16338),
    .O(net_16362)
  );
  Odrv4 odrv_4_12_16454_16487 (
    .I(net_16454),
    .O(net_16487)
  );
  Odrv4 odrv_4_12_16455_16598 (
    .I(net_16455),
    .O(net_16598)
  );
  Odrv4 odrv_4_12_16457_20435 (
    .I(net_16457),
    .O(net_20435)
  );
  Odrv4 odrv_4_12_16458_12758 (
    .I(net_16458),
    .O(net_12758)
  );
  Odrv4 odrv_4_12_16459_16481 (
    .I(net_16459),
    .O(net_16481)
  );
  Odrv4 odrv_4_12_16461_16611 (
    .I(net_16461),
    .O(net_16611)
  );
  Odrv4 odrv_4_13_16584_16717 (
    .I(net_16584),
    .O(net_16717)
  );
  Odrv4 odrv_4_14_16701_20311 (
    .I(net_16701),
    .O(net_20311)
  );
  Odrv4 odrv_4_14_16707_16603 (
    .I(net_16707),
    .O(net_16603)
  );
  Odrv4 odrv_4_17_17069_21035 (
    .I(net_17069),
    .O(net_21035)
  );
  Odrv4 odrv_4_17_17073_21045 (
    .I(net_17073),
    .O(net_21045)
  );
  Odrv4 odrv_4_17_17075_17205 (
    .I(net_17075),
    .O(net_17205)
  );
  Odrv4 odrv_4_17_17076_20930 (
    .I(net_17076),
    .O(net_20930)
  );
  Odrv4 odrv_4_18_17195_16977 (
    .I(net_17195),
    .O(net_16977)
  );
  Odrv4 odrv_4_19_17315_17220 (
    .I(net_17315),
    .O(net_17220)
  );
  Odrv4 odrv_4_19_17322_17218 (
    .I(net_17322),
    .O(net_17218)
  );
  Odrv4 odrv_4_1_15063_15244 (
    .I(net_15063),
    .O(net_15244)
  );
  Odrv4 odrv_4_1_15063_19076 (
    .I(net_15063),
    .O(net_19076)
  );
  Odrv4 odrv_4_1_15064_19079 (
    .I(net_15064),
    .O(net_19079)
  );
  Odrv4 odrv_4_1_15065_19081 (
    .I(net_15065),
    .O(net_19081)
  );
  Odrv4 odrv_4_22_17690_17585 (
    .I(net_17690),
    .O(net_17585)
  );
  Odrv12 odrv_4_31_18791_21280 (
    .I(net_18791),
    .O(net_21280)
  );
  Odrv4 odrv_4_3_15352_7176 (
    .I(net_15352),
    .O(net_7176)
  );
  Odrv4 odrv_4_4_15470_15243 (
    .I(net_15470),
    .O(net_15243)
  );
  Odrv4 odrv_4_4_15471_19440 (
    .I(net_15471),
    .O(net_19440)
  );
  Odrv4 odrv_4_4_15472_19442 (
    .I(net_15472),
    .O(net_19442)
  );
  Odrv4 odrv_4_4_15473_15250 (
    .I(net_15473),
    .O(net_15250)
  );
  Odrv4 odrv_4_4_15473_19080 (
    .I(net_15473),
    .O(net_19080)
  );
  Odrv4 odrv_4_4_15475_11778 (
    .I(net_15475),
    .O(net_11778)
  );
  Odrv4 odrv_4_5_15594_15737 (
    .I(net_15594),
    .O(net_15737)
  );
  Odrv4 odrv_4_5_15595_15739 (
    .I(net_15595),
    .O(net_15739)
  );
  Odrv4 odrv_4_5_15598_15746 (
    .I(net_15598),
    .O(net_15746)
  );
  Odrv4 odrv_4_5_15598_19561 (
    .I(net_15598),
    .O(net_19561)
  );
  Odrv4 odrv_4_5_15599_11903 (
    .I(net_15599),
    .O(net_11903)
  );
  Odrv4 odrv_4_5_15599_15622 (
    .I(net_15599),
    .O(net_15622)
  );
  Odrv4 odrv_4_5_15599_15729 (
    .I(net_15599),
    .O(net_15729)
  );
  Odrv4 odrv_4_5_15599_15748 (
    .I(net_15599),
    .O(net_15748)
  );
  Odrv4 odrv_4_6_15720_19699 (
    .I(net_15720),
    .O(net_19699)
  );
  Odrv4 odrv_4_7_15839_19805 (
    .I(net_15839),
    .O(net_19805)
  );
  Odrv4 odrv_4_7_15841_19811 (
    .I(net_15841),
    .O(net_19811)
  );
  Odrv4 odrv_4_7_15843_19456 (
    .I(net_15843),
    .O(net_19456)
  );
  Odrv4 odrv_4_8_15969_19951 (
    .I(net_15969),
    .O(net_19951)
  );
  Odrv4 odrv_4_9_16085_12399 (
    .I(net_16085),
    .O(net_12399)
  );
  Odrv4 odrv_4_9_16086_19950 (
    .I(net_16086),
    .O(net_19950)
  );
  Odrv4 odrv_4_9_16087_16231 (
    .I(net_16087),
    .O(net_16231)
  );
  Odrv4 odrv_4_9_16088_16223 (
    .I(net_16088),
    .O(net_16223)
  );
  Odrv4 odrv_4_9_16089_12389 (
    .I(net_16089),
    .O(net_12389)
  );
  Odrv4 odrv_4_9_16090_19942 (
    .I(net_16090),
    .O(net_19942)
  );
  Odrv4 odrv_4_9_16091_19944 (
    .I(net_16091),
    .O(net_19944)
  );
  Odrv4 odrv_4_9_16092_16225 (
    .I(net_16092),
    .O(net_16225)
  );
  Odrv4 odrv_5_10_20039_20181 (
    .I(net_20039),
    .O(net_20181)
  );
  Odrv4 odrv_5_10_20040_23778 (
    .I(net_20040),
    .O(net_23778)
  );
  Odrv4 odrv_5_10_20041_19948 (
    .I(net_20041),
    .O(net_19948)
  );
  Odrv4 odrv_5_10_20042_24020 (
    .I(net_20042),
    .O(net_24020)
  );
  Odrv4 odrv_5_10_20043_20190 (
    .I(net_20043),
    .O(net_20190)
  );
  Odrv4 odrv_5_10_20044_24007 (
    .I(net_20044),
    .O(net_24007)
  );
  Odrv12 odrv_5_10_20045_23266 (
    .I(net_20045),
    .O(net_23266)
  );
  Odrv4 odrv_5_10_20046_23774 (
    .I(net_20046),
    .O(net_23774)
  );
  Odrv4 odrv_5_11_20162_16476 (
    .I(net_20162),
    .O(net_16476)
  );
  Odrv4 odrv_5_11_20162_20195 (
    .I(net_20162),
    .O(net_20195)
  );
  Odrv4 odrv_5_11_20163_20306 (
    .I(net_20163),
    .O(net_20306)
  );
  Odrv4 odrv_5_11_20164_19945 (
    .I(net_20164),
    .O(net_19945)
  );
  Odrv4 odrv_5_11_20164_20309 (
    .I(net_20164),
    .O(net_20309)
  );
  Odrv4 odrv_5_11_20165_24136 (
    .I(net_20165),
    .O(net_24136)
  );
  Odrv4 odrv_5_11_20166_20187 (
    .I(net_20166),
    .O(net_20187)
  );
  Odrv4 odrv_5_11_20167_20189 (
    .I(net_20167),
    .O(net_20189)
  );
  Odrv4 odrv_5_11_20168_20191 (
    .I(net_20168),
    .O(net_20191)
  );
  Odrv4 odrv_5_11_20169_20319 (
    .I(net_20169),
    .O(net_20319)
  );
  Odrv4 odrv_5_12_20285_16599 (
    .I(net_20285),
    .O(net_16599)
  );
  Odrv12 odrv_5_12_20285_22746 (
    .I(net_20285),
    .O(net_22746)
  );
  Odrv4 odrv_5_12_20285_24148 (
    .I(net_20285),
    .O(net_24148)
  );
  Odrv4 odrv_5_12_20286_16591 (
    .I(net_20286),
    .O(net_16591)
  );
  Odrv4 odrv_5_12_20286_20066 (
    .I(net_20286),
    .O(net_20066)
  );
  Odrv4 odrv_5_12_20286_20429 (
    .I(net_20286),
    .O(net_20429)
  );
  Odrv4 odrv_5_12_20286_24024 (
    .I(net_20286),
    .O(net_24024)
  );
  Odrv4 odrv_5_12_20288_20070 (
    .I(net_20288),
    .O(net_20070)
  );
  Odrv4 odrv_5_12_20288_20423 (
    .I(net_20288),
    .O(net_20423)
  );
  Odrv4 odrv_5_12_20290_20312 (
    .I(net_20290),
    .O(net_20312)
  );
  Odrv4 odrv_5_12_20291_16595 (
    .I(net_20291),
    .O(net_16595)
  );
  Odrv4 odrv_5_12_20292_12761 (
    .I(net_20292),
    .O(net_12761)
  );
  Odrv4 odrv_5_12_20292_24146 (
    .I(net_20292),
    .O(net_24146)
  );
  Odrv4 odrv_5_13_20408_20313 (
    .I(net_20408),
    .O(net_20313)
  );
  Odrv12 odrv_5_13_20408_22861 (
    .I(net_20408),
    .O(net_22861)
  );
  Odrv4 odrv_5_13_20408_24145 (
    .I(net_20408),
    .O(net_24145)
  );
  Odrv4 odrv_5_13_20409_20443 (
    .I(net_20409),
    .O(net_20443)
  );
  Odrv4 odrv_5_13_20409_20552 (
    .I(net_20409),
    .O(net_20552)
  );
  Odrv4 odrv_5_13_20409_24147 (
    .I(net_20409),
    .O(net_24147)
  );
  Odrv4 odrv_5_13_20410_20317 (
    .I(net_20410),
    .O(net_20317)
  );
  Odrv4 odrv_5_14_20531_24268 (
    .I(net_20531),
    .O(net_24268)
  );
  Odrv4 odrv_5_14_20538_24392 (
    .I(net_20538),
    .O(net_24392)
  );
  Odrv4 odrv_5_15_20656_20437 (
    .I(net_20656),
    .O(net_20437)
  );
  Odrv4 odrv_5_15_20659_24639 (
    .I(net_20659),
    .O(net_24639)
  );
  Odrv4 odrv_5_16_20779_20560 (
    .I(net_20779),
    .O(net_20560)
  );
  Odrv4 odrv_5_16_20782_20566 (
    .I(net_20782),
    .O(net_20566)
  );
  Odrv4 odrv_5_16_20783_20806 (
    .I(net_20783),
    .O(net_20806)
  );
  Odrv4 odrv_5_16_20784_24512 (
    .I(net_20784),
    .O(net_24512)
  );
  Odrv4 odrv_5_17_20901_17206 (
    .I(net_20901),
    .O(net_17206)
  );
  Odrv4 odrv_5_17_20901_24870 (
    .I(net_20901),
    .O(net_24870)
  );
  Odrv4 odrv_5_18_21024_24634 (
    .I(net_21024),
    .O(net_24634)
  );
  Odrv4 odrv_5_18_21026_21161 (
    .I(net_21026),
    .O(net_21161)
  );
  Odrv4 odrv_5_18_21027_17327 (
    .I(net_21027),
    .O(net_17327)
  );
  Odrv4 odrv_5_19_21150_17450 (
    .I(net_21150),
    .O(net_17450)
  );
  Odrv4 odrv_5_2_19020_22898 (
    .I(net_19020),
    .O(net_22898)
  );
  Odrv12 odrv_5_31_22622_25111 (
    .I(net_22622),
    .O(net_25111)
  );
  Odrv4 odrv_5_31_22622_26489 (
    .I(net_22622),
    .O(net_26489)
  );
  Odrv4 odrv_5_3_19182_19069 (
    .I(net_19182),
    .O(net_19069)
  );
  Odrv4 odrv_5_3_19185_19209 (
    .I(net_19185),
    .O(net_19209)
  );
  Odrv4 odrv_5_4_19301_19334 (
    .I(net_19301),
    .O(net_19334)
  );
  Odrv4 odrv_5_4_19302_19336 (
    .I(net_19302),
    .O(net_19336)
  );
  Odrv4 odrv_5_4_19303_19448 (
    .I(net_19303),
    .O(net_19448)
  );
  Odrv4 odrv_5_4_19303_23273 (
    .I(net_19303),
    .O(net_23273)
  );
  Odrv4 odrv_5_4_19304_19450 (
    .I(net_19304),
    .O(net_19450)
  );
  Odrv4 odrv_5_4_19305_19326 (
    .I(net_19305),
    .O(net_19326)
  );
  Odrv4 odrv_5_4_19306_23286 (
    .I(net_19306),
    .O(net_23286)
  );
  Odrv4 odrv_5_4_19307_23288 (
    .I(net_19307),
    .O(net_23288)
  );
  Odrv4 odrv_5_4_19308_19441 (
    .I(net_19308),
    .O(net_19441)
  );
  Odrv4 odrv_5_5_19425_15730 (
    .I(net_19425),
    .O(net_15730)
  );
  Odrv4 odrv_5_5_19426_11898 (
    .I(net_19426),
    .O(net_11898)
  );
  Odrv4 odrv_5_5_19427_11902 (
    .I(net_19427),
    .O(net_11902)
  );
  Odrv4 odrv_5_5_19428_11904 (
    .I(net_19428),
    .O(net_11904)
  );
  Odrv4 odrv_5_5_19429_23392 (
    .I(net_19429),
    .O(net_23392)
  );
  Odrv4 odrv_5_5_19430_23157 (
    .I(net_19430),
    .O(net_23157)
  );
  Odrv4 odrv_5_6_19554_15859 (
    .I(net_19554),
    .O(net_15859)
  );
  Odrv4 odrv_5_7_19671_19814 (
    .I(net_19671),
    .O(net_19814)
  );
  Odrv12 odrv_5_7_19672_23389 (
    .I(net_19672),
    .O(net_23389)
  );
  Odrv4 odrv_5_7_19675_23289 (
    .I(net_19675),
    .O(net_23289)
  );
  Odrv4 odrv_5_8_19793_23402 (
    .I(net_19793),
    .O(net_23402)
  );
  Odrv4 odrv_5_8_19794_19574 (
    .I(net_19794),
    .O(net_19574)
  );
  Odrv4 odrv_5_8_19795_19939 (
    .I(net_19795),
    .O(net_19939)
  );
  Odrv4 odrv_5_8_19796_23536 (
    .I(net_19796),
    .O(net_23536)
  );
  Odrv4 odrv_5_8_19796_23767 (
    .I(net_19796),
    .O(net_23767)
  );
  Odrv4 odrv_5_8_19797_23769 (
    .I(net_19797),
    .O(net_23769)
  );
  Odrv4 odrv_5_8_19800_19933 (
    .I(net_19800),
    .O(net_19933)
  );
  Odrv4 odrv_5_9_19916_20058 (
    .I(net_19916),
    .O(net_20058)
  );
  Odrv4 odrv_5_9_19916_23779 (
    .I(net_19916),
    .O(net_23779)
  );
  Odrv12 odrv_5_9_19917_1991 (
    .I(net_19917),
    .O(net_1991)
  );
  Odrv4 odrv_5_9_19917_23781 (
    .I(net_19917),
    .O(net_23781)
  );
  Odrv4 odrv_5_9_19918_20062 (
    .I(net_19918),
    .O(net_20062)
  );
  Odrv4 odrv_5_9_19918_20063 (
    .I(net_19918),
    .O(net_20063)
  );
  Odrv4 odrv_5_9_19919_20054 (
    .I(net_19919),
    .O(net_20054)
  );
  Odrv4 odrv_5_9_19919_20065 (
    .I(net_19919),
    .O(net_20065)
  );
  Odrv4 odrv_5_9_19920_20067 (
    .I(net_19920),
    .O(net_20067)
  );
  Odrv4 odrv_5_9_19920_23771 (
    .I(net_19920),
    .O(net_23771)
  );
  Odrv4 odrv_5_9_19921_20069 (
    .I(net_19921),
    .O(net_20069)
  );
  Odrv4 odrv_5_9_19921_23773 (
    .I(net_19921),
    .O(net_23773)
  );
  Odrv4 odrv_5_9_19922_20071 (
    .I(net_19922),
    .O(net_20071)
  );
  Odrv4 odrv_5_9_19922_23775 (
    .I(net_19922),
    .O(net_23775)
  );
  Odrv4 odrv_5_9_19923_20073 (
    .I(net_19923),
    .O(net_20073)
  );
  Odrv4 odrv_6_0_22846_18923 (
    .I(net_22846),
    .O(net_18923)
  );
  Odrv4 odrv_6_0_22846_22874 (
    .I(net_22846),
    .O(net_22874)
  );
  Odrv4 odrv_6_0_22848_22756 (
    .I(net_22848),
    .O(net_22756)
  );
  Odrv4 odrv_6_0_22848_22895 (
    .I(net_22848),
    .O(net_22895)
  );
  Odrv4 odrv_6_10_23874_27635 (
    .I(net_23874),
    .O(net_27635)
  );
  Odrv4 odrv_6_10_23875_27627 (
    .I(net_23875),
    .O(net_27627)
  );
  Odrv4 odrv_6_10_23876_24006 (
    .I(net_23876),
    .O(net_24006)
  );
  Odrv4 odrv_6_11_23994_27731 (
    .I(net_23994),
    .O(net_27731)
  );
  Odrv4 odrv_6_11_23996_16471 (
    .I(net_23996),
    .O(net_16471)
  );
  Odrv4 odrv_6_11_23999_16477 (
    .I(net_23999),
    .O(net_16477)
  );
  Odrv4 odrv_6_11_24000_16469 (
    .I(net_24000),
    .O(net_16469)
  );
  Odrv4 odrv_6_12_24117_20422 (
    .I(net_24117),
    .O(net_20422)
  );
  Odrv4 odrv_6_12_24118_24263 (
    .I(net_24118),
    .O(net_24263)
  );
  Odrv4 odrv_6_12_24119_24265 (
    .I(net_24119),
    .O(net_24265)
  );
  Odrv4 odrv_6_12_24121_23905 (
    .I(net_24121),
    .O(net_23905)
  );
  Odrv4 odrv_6_12_24122_20426 (
    .I(net_24122),
    .O(net_20426)
  );
  Odrv4 odrv_6_12_24123_24256 (
    .I(net_24123),
    .O(net_24256)
  );
  Odrv4 odrv_6_31_26453_26358 (
    .I(net_26453),
    .O(net_26358)
  );
  Odrv12 odrv_6_31_26453_28542 (
    .I(net_26453),
    .O(net_28542)
  );
  Odrv4 odrv_6_31_26453_29689 (
    .I(net_26453),
    .O(net_29689)
  );
  Odrv4 odrv_6_4_23134_15606 (
    .I(net_23134),
    .O(net_15606)
  );
  Odrv4 odrv_6_4_23135_27028 (
    .I(net_23135),
    .O(net_27028)
  );
  Odrv4 odrv_6_4_23136_23283 (
    .I(net_23136),
    .O(net_23283)
  );
  Odrv4 odrv_6_4_23137_27032 (
    .I(net_23137),
    .O(net_27032)
  );
  Odrv4 odrv_6_4_23138_23287 (
    .I(net_23138),
    .O(net_23287)
  );
  Odrv4 odrv_6_4_23139_15608 (
    .I(net_23139),
    .O(net_15608)
  );
  Odrv4 odrv_6_9_23748_23782 (
    .I(net_23748),
    .O(net_23782)
  );
  Odrv12 odrv_6_9_23750_2002 (
    .I(net_23750),
    .O(net_2002)
  );
  Odrv4 odrv_6_9_23751_16227 (
    .I(net_23751),
    .O(net_16227)
  );
  Odrv12 odrv_6_9_23753_2012 (
    .I(net_23753),
    .O(net_2012)
  );
  Odrv12 odrv_6_9_23754_1992 (
    .I(net_23754),
    .O(net_1992)
  );
  Odrv4 odrv_7_10_27484_27338 (
    .I(net_27484),
    .O(net_27338)
  );
  Odrv4 odrv_7_10_27488_27647 (
    .I(net_27488),
    .O(net_27647)
  );
  Odrv4 odrv_7_11_27587_27743 (
    .I(net_27587),
    .O(net_27743)
  );
  Odrv4 odrv_7_11_27588_27640 (
    .I(net_27588),
    .O(net_27640)
  );
  Odrv4 odrv_7_13_27790_31054 (
    .I(net_27790),
    .O(net_31054)
  );
  Odrv4 odrv_7_13_27793_27739 (
    .I(net_27793),
    .O(net_27739)
  );
  Odrv4 odrv_7_13_27793_31172 (
    .I(net_27793),
    .O(net_31172)
  );
  Odrv4 odrv_7_14_27892_27746 (
    .I(net_27892),
    .O(net_27746)
  );
  Odrv4 odrv_7_14_27892_28036 (
    .I(net_27892),
    .O(net_28036)
  );
  Odrv4 odrv_7_14_27892_31177 (
    .I(net_27892),
    .O(net_31177)
  );
  Odrv4 odrv_7_14_27893_31179 (
    .I(net_27893),
    .O(net_31179)
  );
  Odrv4 odrv_7_15_27991_27947 (
    .I(net_27991),
    .O(net_27947)
  );
  Odrv4 odrv_7_15_27992_27844 (
    .I(net_27992),
    .O(net_27844)
  );
  Odrv4 odrv_7_15_27994_31300 (
    .I(net_27994),
    .O(net_31300)
  );
  Odrv4 odrv_7_15_27995_27850 (
    .I(net_27995),
    .O(net_27850)
  );
  Odrv4 odrv_7_15_27996_31304 (
    .I(net_27996),
    .O(net_31304)
  );
  Odrv4 odrv_7_15_27997_27943 (
    .I(net_27997),
    .O(net_27943)
  );
  Odrv4 odrv_7_15_27998_31546 (
    .I(net_27998),
    .O(net_31546)
  );
  Odrv4 odrv_7_17_28202_21038 (
    .I(net_28202),
    .O(net_21038)
  );
  Odrv4 odrv_7_3_26767_30175 (
    .I(net_26767),
    .O(net_30175)
  );
  Odrv4 odrv_7_3_26770_26914 (
    .I(net_26770),
    .O(net_26914)
  );
  Odrv4 odrv_7_3_26771_30185 (
    .I(net_26771),
    .O(net_30185)
  );
  Odrv4 odrv_7_4_26872_26721 (
    .I(net_26872),
    .O(net_26721)
  );
  Odrv4 odrv_7_4_26874_19445 (
    .I(net_26874),
    .O(net_19445)
  );
  Odrv4 odrv_7_4_26874_30189 (
    .I(net_26874),
    .O(net_30189)
  );
  Odrv4 odrv_7_4_26876_30321 (
    .I(net_26876),
    .O(net_30321)
  );
  Odrv4 odrv_7_5_26975_23390 (
    .I(net_26975),
    .O(net_23390)
  );
  Odrv4 odrv_7_5_26975_30310 (
    .I(net_26975),
    .O(net_30310)
  );
  Odrv4 odrv_7_5_26977_27135 (
    .I(net_26977),
    .O(net_27135)
  );
  Odrv4 odrv_7_6_27074_23515 (
    .I(net_27074),
    .O(net_23515)
  );
  Odrv4 odrv_7_6_27077_19689 (
    .I(net_27077),
    .O(net_19689)
  );
  Odrv4 odrv_7_6_27078_23517 (
    .I(net_27078),
    .O(net_23517)
  );
  Odrv4 odrv_7_6_27078_27235 (
    .I(net_27078),
    .O(net_27235)
  );
  Odrv4 odrv_7_6_27079_19693 (
    .I(net_27079),
    .O(net_19693)
  );
  Odrv4 odrv_7_6_27079_27025 (
    .I(net_27079),
    .O(net_27025)
  );
  Odrv4 odrv_7_7_27179_23636 (
    .I(net_27179),
    .O(net_23636)
  );
  Odrv4 odrv_7_7_27180_23640 (
    .I(net_27180),
    .O(net_23640)
  );
  Odrv4 odrv_7_8_27280_27435 (
    .I(net_27280),
    .O(net_27435)
  );
  Odrv12 odrv_7_9_27379_30420 (
    .I(net_27379),
    .O(net_30420)
  );
  Odrv4 odrv_7_9_27380_27444 (
    .I(net_27380),
    .O(net_27444)
  );
  Odrv4 odrv_7_9_27381_27535 (
    .I(net_27381),
    .O(net_27535)
  );
  Odrv4 odrv_7_9_27382_27537 (
    .I(net_27382),
    .O(net_27537)
  );
  Odrv4 odrv_7_9_27383_23882 (
    .I(net_27383),
    .O(net_23882)
  );
  Odrv4 odrv_7_9_27385_27524 (
    .I(net_27385),
    .O(net_27524)
  );
  Odrv12 odrv_7_9_27386_30296 (
    .I(net_27386),
    .O(net_30296)
  );
  Odrv4 odrv_8_10_30902_30936 (
    .I(net_30902),
    .O(net_30936)
  );
  Odrv4 odrv_8_10_30903_31048 (
    .I(net_30903),
    .O(net_31048)
  );
  Odrv4 odrv_8_11_31029_30813 (
    .I(net_31029),
    .O(net_30813)
  );
  Odrv4 odrv_8_11_31031_30927 (
    .I(net_31031),
    .O(net_30927)
  );
  Odrv4 odrv_8_11_31031_31164 (
    .I(net_31031),
    .O(net_31164)
  );
  Odrv4 odrv_8_11_31031_34759 (
    .I(net_31031),
    .O(net_34759)
  );
  Odrv4 odrv_8_12_31154_34882 (
    .I(net_31154),
    .O(net_34882)
  );
  Odrv4 odrv_8_13_31271_31051 (
    .I(net_31271),
    .O(net_31051)
  );
  Odrv4 odrv_8_13_31272_31053 (
    .I(net_31272),
    .O(net_31053)
  );
  Odrv4 odrv_8_13_31277_35131 (
    .I(net_31277),
    .O(net_35131)
  );
  Odrv4 odrv_8_15_31516_35482 (
    .I(net_31516),
    .O(net_35482)
  );
  Odrv4 odrv_8_15_31517_35127 (
    .I(net_31517),
    .O(net_35127)
  );
  Odrv4 odrv_8_15_31518_35488 (
    .I(net_31518),
    .O(net_35488)
  );
  Odrv4 odrv_8_15_31519_35497 (
    .I(net_31519),
    .O(net_35497)
  );
  Odrv4 odrv_8_15_31520_35499 (
    .I(net_31520),
    .O(net_35499)
  );
  Odrv4 odrv_8_15_31522_31652 (
    .I(net_31522),
    .O(net_31652)
  );
  Odrv4 odrv_8_15_31523_35251 (
    .I(net_31523),
    .O(net_35251)
  );
  Odrv4 odrv_8_16_31640_35378 (
    .I(net_31640),
    .O(net_35378)
  );
  Odrv4 odrv_8_16_31642_35254 (
    .I(net_31642),
    .O(net_35254)
  );
  Odrv4 odrv_8_16_31645_35372 (
    .I(net_31645),
    .O(net_35372)
  );
  Odrv4 odrv_8_2_29883_33889 (
    .I(net_29883),
    .O(net_33889)
  );
  Odrv4 odrv_8_2_29887_33771 (
    .I(net_29887),
    .O(net_33771)
  );
  Odrv12 odrv_8_31_33484_35973 (
    .I(net_33484),
    .O(net_35973)
  );
  Odrv12 odrv_8_31_33486_36219 (
    .I(net_33486),
    .O(net_36219)
  );
  Odrv4 odrv_8_3_30040_30182 (
    .I(net_30040),
    .O(net_30182)
  );
  Odrv4 odrv_8_3_30046_30069 (
    .I(net_30046),
    .O(net_30069)
  );
  Odrv4 odrv_8_4_30163_30305 (
    .I(net_30163),
    .O(net_30305)
  );
  Odrv4 odrv_8_4_30166_30301 (
    .I(net_30166),
    .O(net_30301)
  );
  Odrv4 odrv_8_4_30169_33896 (
    .I(net_30169),
    .O(net_33896)
  );
  Odrv4 odrv_8_4_30170_34152 (
    .I(net_30170),
    .O(net_34152)
  );
  Odrv4 odrv_8_5_30286_34252 (
    .I(net_30286),
    .O(net_34252)
  );
  Odrv4 odrv_8_5_30288_23391 (
    .I(net_30288),
    .O(net_23391)
  );
  Odrv12 odrv_8_5_30292_33605 (
    .I(net_30292),
    .O(net_33605)
  );
  Odrv4 odrv_8_6_30409_30442 (
    .I(net_30409),
    .O(net_30442)
  );
  Odrv4 odrv_8_6_30410_34148 (
    .I(net_30410),
    .O(net_34148)
  );
  Odrv4 odrv_8_6_30412_30320 (
    .I(net_30412),
    .O(net_30320)
  );
  Odrv4 odrv_8_6_30413_30560 (
    .I(net_30413),
    .O(net_30560)
  );
  Odrv4 odrv_8_6_30414_30436 (
    .I(net_30414),
    .O(net_30436)
  );
  Odrv4 odrv_8_6_30415_30564 (
    .I(net_30415),
    .O(net_30564)
  );
  Odrv4 odrv_8_6_30416_30440 (
    .I(net_30416),
    .O(net_30440)
  );
  Odrv4 odrv_8_7_30532_30565 (
    .I(net_30532),
    .O(net_30565)
  );
  Odrv12 odrv_8_7_30534_34251 (
    .I(net_30534),
    .O(net_34251)
  );
  Odrv4 odrv_8_7_30538_34391 (
    .I(net_30538),
    .O(net_34391)
  );
  Odrv4 odrv_8_9_30778_34387 (
    .I(net_30778),
    .O(net_34387)
  );
  Odrv4 odrv_9_10_34732_34511 (
    .I(net_34732),
    .O(net_34511)
  );
  Odrv4 odrv_9_10_34739_34889 (
    .I(net_34739),
    .O(net_34889)
  );
  Odrv4 odrv_9_10_34739_38593 (
    .I(net_34739),
    .O(net_38593)
  );
  Odrv4 odrv_9_11_34855_31169 (
    .I(net_34855),
    .O(net_31169)
  );
  Odrv4 odrv_9_11_34855_34634 (
    .I(net_34855),
    .O(net_34634)
  );
  Odrv4 odrv_9_11_34855_34760 (
    .I(net_34855),
    .O(net_34760)
  );
  Odrv4 odrv_9_11_34855_34997 (
    .I(net_34855),
    .O(net_34997)
  );
  Odrv4 odrv_9_11_34855_38464 (
    .I(net_34855),
    .O(net_38464)
  );
  Odrv4 odrv_9_11_34855_38592 (
    .I(net_34855),
    .O(net_38592)
  );
  Odrv4 odrv_9_11_34861_27738 (
    .I(net_34861),
    .O(net_27738)
  );
  Odrv4 odrv_9_11_34861_31165 (
    .I(net_34861),
    .O(net_31165)
  );
  Odrv4 odrv_9_11_34861_34756 (
    .I(net_34861),
    .O(net_34756)
  );
  Odrv4 odrv_9_11_34861_34884 (
    .I(net_34861),
    .O(net_34884)
  );
  Odrv4 odrv_9_11_34861_34991 (
    .I(net_34861),
    .O(net_34991)
  );
  Odrv4 odrv_9_11_34861_35010 (
    .I(net_34861),
    .O(net_35010)
  );
  Odrv4 odrv_9_11_34861_38588 (
    .I(net_34861),
    .O(net_38588)
  );
  Odrv4 odrv_9_12_34978_35120 (
    .I(net_34978),
    .O(net_35120)
  );
  Odrv4 odrv_9_12_34979_35122 (
    .I(net_34979),
    .O(net_35122)
  );
  Odrv4 odrv_9_12_34982_35129 (
    .I(net_34982),
    .O(net_35129)
  );
  Odrv4 odrv_9_13_35106_39069 (
    .I(net_35106),
    .O(net_39069)
  );
  Odrv4 odrv_9_13_35107_35130 (
    .I(net_35107),
    .O(net_35130)
  );
  Odrv4 odrv_9_14_35229_31532 (
    .I(net_35229),
    .O(net_31532)
  );
  Odrv4 odrv_9_15_35349_28136 (
    .I(net_35349),
    .O(net_28136)
  );
  Odrv4 odrv_9_16_35470_39436 (
    .I(net_35470),
    .O(net_39436)
  );
  Odrv4 odrv_9_16_35473_35619 (
    .I(net_35473),
    .O(net_35619)
  );
  Odrv4 odrv_9_16_35474_39453 (
    .I(net_35474),
    .O(net_39453)
  );
  Odrv4 odrv_9_16_35475_39455 (
    .I(net_35475),
    .O(net_39455)
  );
  Odrv4 odrv_9_16_35477_39331 (
    .I(net_35477),
    .O(net_39331)
  );
  Odrv4 odrv_9_17_35594_39458 (
    .I(net_35594),
    .O(net_39458)
  );
  Odrv4 odrv_9_18_35717_39581 (
    .I(net_35717),
    .O(net_39581)
  );
  Odrv4 odrv_9_3_33877_33900 (
    .I(net_33877),
    .O(net_33900)
  );
  Odrv4 odrv_9_4_33994_30308 (
    .I(net_33994),
    .O(net_30308)
  );
  Odrv4 odrv_9_4_33999_30302 (
    .I(net_33999),
    .O(net_30302)
  );
  Odrv4 odrv_9_5_34118_30423 (
    .I(net_34118),
    .O(net_30423)
  );
  Odrv4 odrv_9_5_34121_33904 (
    .I(net_34121),
    .O(net_33904)
  );
  Odrv4 odrv_9_5_34124_27118 (
    .I(net_34124),
    .O(net_27118)
  );
  Odrv4 odrv_9_6_34243_34378 (
    .I(net_34243),
    .O(net_34378)
  );
  Odrv4 odrv_9_6_34244_37857 (
    .I(net_34244),
    .O(net_37857)
  );
  Odrv4 odrv_9_7_34364_34507 (
    .I(net_34364),
    .O(net_34507)
  );
  Odrv4 odrv_9_7_34364_37974 (
    .I(net_34364),
    .O(net_37974)
  );
  Odrv4 odrv_9_7_34364_38228 (
    .I(net_34364),
    .O(net_38228)
  );
  Odrv12 odrv_9_7_34368_1555 (
    .I(net_34368),
    .O(net_1555)
  );
  Odrv12 odrv_9_7_34368_37438 (
    .I(net_34368),
    .O(net_37438)
  );
  Odrv4 odrv_9_8_34493_30798 (
    .I(net_34493),
    .O(net_30798)
  );
  Odrv4 odrv_9_8_34493_34389 (
    .I(net_34493),
    .O(net_34389)
  );
  Odrv4 odrv_9_9_34615_34510 (
    .I(net_34615),
    .O(net_34510)
  );
  Odrv4 odrv_9_9_34616_34640 (
    .I(net_34616),
    .O(net_34640)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_12_31_1 (
    .CLOCKENABLE(),
    .DIN0(net_48810),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_12_31_1_dout),
    .PADOEN(io_pad_12_31_1_oe),
    .PADOUT(io_pad_12_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_13_0_1 (
    .CLOCKENABLE(),
    .DIN0(net_49034),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_13_0_1_dout),
    .PADOEN(io_pad_13_0_1_oe),
    .PADOUT(io_pad_13_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_13_31_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_56515),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_13_31_0_dout),
    .PADOEN(io_pad_13_31_0_oe),
    .PADOUT(io_pad_13_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_13_31_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_56518),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_13_31_1_dout),
    .PADOEN(io_pad_13_31_1_oe),
    .PADOUT(io_pad_13_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_15_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_56693),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_15_0_0_dout),
    .PADOEN(io_pad_15_0_0_oe),
    .PADOUT(io_pad_15_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_16_0_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_64205),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_16_0_0_dout),
    .PADOEN(io_pad_16_0_0_oe),
    .PADOUT(io_pad_16_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_16_31_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_68006),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_16_31_0_dout),
    .PADOEN(io_pad_16_31_0_oe),
    .PADOUT(io_pad_16_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_16_31_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_68009),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_16_31_1_dout),
    .PADOEN(io_pad_16_31_1_oe),
    .PADOUT(io_pad_16_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_17_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_64354),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_17_0_0_dout),
    .PADOEN(io_pad_17_0_0_oe),
    .PADOUT(io_pad_17_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_17_31_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_71837),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_17_31_0_dout),
    .PADOEN(io_pad_17_31_0_oe),
    .PADOUT(io_pad_17_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_18_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_68185),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_0_0_dout),
    .PADOEN(io_pad_18_0_0_oe),
    .PADOUT(io_pad_18_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_18_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_71870),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_0_1_dout),
    .PADOEN(io_pad_18_0_1_oe),
    .PADOUT(io_pad_18_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_18_31_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_75668),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_31_0_dout),
    .PADOEN(io_pad_18_31_0_oe),
    .PADOUT(io_pad_18_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_18_31_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_75671),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_31_1_dout),
    .PADOEN(io_pad_18_31_1_oe),
    .PADOUT(io_pad_18_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_19_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_72016),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_19_0_0_dout),
    .PADOEN(io_pad_19_0_0_oe),
    .PADOUT(io_pad_19_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_19_0_1 (
    .CLOCKENABLE(),
    .DIN0(net_72018),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_19_0_1_dout),
    .PADOEN(io_pad_19_0_1_oe),
    .PADOUT(io_pad_19_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_21_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_82732),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_21_0_1_dout),
    .PADOEN(io_pad_21_0_1_oe),
    .PADOUT(io_pad_21_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_22_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_86563),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_22_0_1_dout),
    .PADOEN(io_pad_22_0_1_oe),
    .PADOUT(io_pad_22_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_23_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_86709),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_23_0_0_dout),
    .PADOEN(io_pad_23_0_0_oe),
    .PADOUT(io_pad_23_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_23_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_90394),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_23_0_1_dout),
    .PADOEN(io_pad_23_0_1_oe),
    .PADOUT(io_pad_23_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_4_31_0 (
    .CLOCKENABLE(),
    .DIN0(net_18791),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_4_31_0_dout),
    .PADOEN(io_pad_4_31_0_oe),
    .PADOUT(io_pad_4_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_5_0_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_22697),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_5_0_0_dout),
    .PADOEN(io_pad_5_0_0_oe),
    .PADOUT(io_pad_5_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_5_31_0 (
    .CLOCKENABLE(),
    .DIN0(net_22622),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_5_31_0_dout),
    .PADOEN(io_pad_5_31_0_oe),
    .PADOUT(io_pad_5_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_6_0_0 (
    .CLOCKENABLE(),
    .DIN0(net_22846),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_6_0_0_dout),
    .PADOEN(io_pad_6_0_0_oe),
    .PADOUT(io_pad_6_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_6_0_1 (
    .CLOCKENABLE(),
    .DIN0(net_22848),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_6_0_1_dout),
    .PADOEN(io_pad_6_0_1_oe),
    .PADOUT(io_pad_6_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_6_31_0 (
    .CLOCKENABLE(),
    .DIN0(net_26453),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_6_31_0_dout),
    .PADOEN(io_pad_6_31_0_oe),
    .PADOUT(io_pad_6_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_7_0_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_29728),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_7_0_0_dout),
    .PADOEN(io_pad_7_0_0_oe),
    .PADOUT(io_pad_7_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_8_0_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_33559),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_8_0_0_dout),
    .PADOEN(io_pad_8_0_0_oe),
    .PADOUT(io_pad_8_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_8_31_0 (
    .CLOCKENABLE(),
    .DIN0(net_33484),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_8_31_0_dout),
    .PADOEN(io_pad_8_31_0_oe),
    .PADOUT(io_pad_8_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_8_31_1 (
    .CLOCKENABLE(),
    .DIN0(net_33486),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_8_31_1_dout),
    .PADOEN(io_pad_8_31_1_oe),
    .PADOUT(io_pad_8_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_9_0_0 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_37390),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_9_0_0_dout),
    .PADOEN(io_pad_9_0_0_oe),
    .PADOUT(io_pad_9_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_9_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_37393),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_9_0_1_dout),
    .PADOEN(io_pad_9_0_1_oe),
    .PADOUT(io_pad_9_0_1_din)
  );
  SB_RAM40_4K ram_6_11 (
    .RCLK(net_27712),
    .RCLKE(net_27713),
    .RE(net_27714),
    .WCLK(net_27814),
    .WCLKE(net_27815),
    .WE(),
    .MASK({dangling_wire_10, dangling_wire_9, dangling_wire_8, dangling_wire_7, dangling_wire_6, dangling_wire_5, dangling_wire_19, dangling_wire_18, dangling_wire_17, dangling_wire_16, dangling_wire_15, dangling_wire_14, dangling_wire_13, dangling_wire_12, dangling_wire_11, dangling_wire_4}),
    .RADDR({dangling_wire_20, dangling_wire_28, dangling_wire_27, dangling_wire_26, dangling_wire_25, dangling_wire_24, dangling_wire_23, dangling_wire_22, dangling_wire_21, net_27702_cascademuxed, net_27701_cascademuxed}),
    .RDATA({net_23993, net_23994, net_23995, net_23996, net_23997, net_23998, net_23999, net_24000, net_24116, net_24117, net_24118, net_24119, net_24120, net_24121, net_24122, net_24123}),
    .WADDR({dangling_wire_30, dangling_wire_39, dangling_wire_38, dangling_wire_37, dangling_wire_36, dangling_wire_35, dangling_wire_34, dangling_wire_33, dangling_wire_32, dangling_wire_31, dangling_wire_29}),
    .WDATA({dangling_wire_46, dangling_wire_45, dangling_wire_44, dangling_wire_43, dangling_wire_42, dangling_wire_41, dangling_wire_55, dangling_wire_54, dangling_wire_53, dangling_wire_52, dangling_wire_51, dangling_wire_50, dangling_wire_49, dangling_wire_48, dangling_wire_47, dangling_wire_40})
  );
  SB_RAM40_4K ram_6_3 (
    .RCLK(net_26896),
    .RCLKE(net_26897),
    .RE(net_26898),
    .WCLK(net_26998),
    .WCLKE(net_26999),
    .WE(net_27008),
    .MASK({net_26882, net_26881, net_26880, net_26879, net_26878, net_26877, net_26884, net_26883, net_26986, net_26985, net_26984, net_26983, net_26982, net_26981, net_26980, net_26979}),
    .RADDR({dangling_wire_56, dangling_wire_60, dangling_wire_59, dangling_wire_58, dangling_wire_57, net_26891_cascademuxed, net_26890_cascademuxed, net_26889_cascademuxed, net_26888_cascademuxed, net_26886_cascademuxed, net_26885_cascademuxed}),
    .RDATA({dangling_wire_64, dangling_wire_63, dangling_wire_62, dangling_wire_61, net_23013, net_23014, net_23015, net_23016, net_23132, net_23133, net_23134, net_23135, net_23136, net_23137, net_23138, net_23139}),
    .WADDR({dangling_wire_65, dangling_wire_69, dangling_wire_68, dangling_wire_67, dangling_wire_66, net_26993_cascademuxed, net_26992_cascademuxed, net_26991_cascademuxed, net_26990_cascademuxed, net_26988_cascademuxed, net_26987_cascademuxed}),
    .WDATA({dangling_wire_73, dangling_wire_72, dangling_wire_71, dangling_wire_70, net_26900, net_26899, net_26906, net_26905, net_27007, net_27006, net_27005, net_27004, net_27003, net_27002, net_27001, net_27000})
  );
  SB_RAM40_4K ram_6_9 (
    .RCLK(net_27508),
    .RCLKE(net_27509),
    .RE(net_27510),
    .WCLK(net_27610),
    .WCLKE(net_27611),
    .WE(),
    .MASK({dangling_wire_80, dangling_wire_79, dangling_wire_78, dangling_wire_77, dangling_wire_76, dangling_wire_75, dangling_wire_89, dangling_wire_88, dangling_wire_87, dangling_wire_86, dangling_wire_85, dangling_wire_84, dangling_wire_83, dangling_wire_82, dangling_wire_81, dangling_wire_74}),
    .RADDR({dangling_wire_90, dangling_wire_98, dangling_wire_97, dangling_wire_96, dangling_wire_95, dangling_wire_94, dangling_wire_93, dangling_wire_92, dangling_wire_91, net_27498_cascademuxed, net_27497_cascademuxed}),
    .RDATA({net_23747, net_23748, net_23749, net_23750, net_23751, net_23752, net_23753, net_23754, net_23870, net_23871, net_23872, net_23873, net_23874, net_23875, net_23876, net_23877}),
    .WADDR({dangling_wire_100, dangling_wire_109, dangling_wire_108, dangling_wire_107, dangling_wire_106, dangling_wire_105, dangling_wire_104, dangling_wire_103, dangling_wire_102, dangling_wire_101, dangling_wire_99}),
    .WDATA({dangling_wire_116, dangling_wire_115, dangling_wire_114, dangling_wire_113, dangling_wire_112, dangling_wire_111, dangling_wire_125, dangling_wire_124, dangling_wire_123, dangling_wire_122, dangling_wire_121, dangling_wire_120, dangling_wire_119, dangling_wire_118, dangling_wire_117, dangling_wire_110})
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t1 (
    .carryinitin(),
    .carryinitout(t0)
  );
  CascadeMux t10 (
    .I(net_6955),
    .O(net_6955_cascademuxed)
  );
  CascadeMux t100 (
    .I(net_12588),
    .O(net_12588_cascademuxed)
  );
  CascadeMux t1000 (
    .I(net_69672),
    .O(net_69672_cascademuxed)
  );
  CascadeMux t1001 (
    .I(net_69678),
    .O(net_69678_cascademuxed)
  );
  CascadeMux t1002 (
    .I(net_69684),
    .O(net_69684_cascademuxed)
  );
  CascadeMux t1003 (
    .I(net_69690),
    .O(net_69690_cascademuxed)
  );
  CascadeMux t1005 (
    .I(net_69696),
    .O(net_69696_cascademuxed)
  );
  CascadeMux t1006 (
    .I(net_69777),
    .O(net_69777_cascademuxed)
  );
  CascadeMux t1007 (
    .I(net_69783),
    .O(net_69783_cascademuxed)
  );
  CascadeMux t1008 (
    .I(net_69789),
    .O(net_69789_cascademuxed)
  );
  CascadeMux t1009 (
    .I(net_69795),
    .O(net_69795_cascademuxed)
  );
  CascadeMux t101 (
    .I(net_12594),
    .O(net_12594_cascademuxed)
  );
  CascadeMux t1010 (
    .I(net_69801),
    .O(net_69801_cascademuxed)
  );
  CascadeMux t1011 (
    .I(net_69813),
    .O(net_69813_cascademuxed)
  );
  CascadeMux t1012 (
    .I(net_69819),
    .O(net_69819_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t1014 (
    .carryinitin(),
    .carryinitout(t1013)
  );
  CascadeMux t1015 (
    .I(net_69900),
    .O(net_69900_cascademuxed)
  );
  CascadeMux t1016 (
    .I(net_69918),
    .O(net_69918_cascademuxed)
  );
  CascadeMux t1017 (
    .I(net_69930),
    .O(net_69930_cascademuxed)
  );
  CascadeMux t1018 (
    .I(net_70023),
    .O(net_70023_cascademuxed)
  );
  CascadeMux t1019 (
    .I(net_70035),
    .O(net_70035_cascademuxed)
  );
  CascadeMux t102 (
    .I(net_12600),
    .O(net_12600_cascademuxed)
  );
  CascadeMux t1020 (
    .I(net_70041),
    .O(net_70041_cascademuxed)
  );
  CascadeMux t1021 (
    .I(net_70152),
    .O(net_70152_cascademuxed)
  );
  CascadeMux t1022 (
    .I(net_70170),
    .O(net_70170_cascademuxed)
  );
  CascadeMux t1023 (
    .I(net_70182),
    .O(net_70182_cascademuxed)
  );
  CascadeMux t1024 (
    .I(net_70188),
    .O(net_70188_cascademuxed)
  );
  CascadeMux t1025 (
    .I(net_72261),
    .O(net_72261_cascademuxed)
  );
  CascadeMux t1026 (
    .I(net_72267),
    .O(net_72267_cascademuxed)
  );
  CascadeMux t1027 (
    .I(net_72279),
    .O(net_72279_cascademuxed)
  );
  CascadeMux t1028 (
    .I(net_72285),
    .O(net_72285_cascademuxed)
  );
  CascadeMux t1029 (
    .I(net_72378),
    .O(net_72378_cascademuxed)
  );
  CascadeMux t103 (
    .I(net_12606),
    .O(net_12606_cascademuxed)
  );
  CascadeMux t1030 (
    .I(net_72384),
    .O(net_72384_cascademuxed)
  );
  CascadeMux t1031 (
    .I(net_72390),
    .O(net_72390_cascademuxed)
  );
  CascadeMux t1032 (
    .I(net_72396),
    .O(net_72396_cascademuxed)
  );
  CascadeMux t1033 (
    .I(net_72402),
    .O(net_72402_cascademuxed)
  );
  CascadeMux t1034 (
    .I(net_72408),
    .O(net_72408_cascademuxed)
  );
  CascadeMux t1035 (
    .I(net_72414),
    .O(net_72414_cascademuxed)
  );
  CascadeMux t1036 (
    .I(net_72420),
    .O(net_72420_cascademuxed)
  );
  CascadeMux t1037 (
    .I(net_72501),
    .O(net_72501_cascademuxed)
  );
  CascadeMux t1038 (
    .I(net_72537),
    .O(net_72537_cascademuxed)
  );
  CascadeMux t1039 (
    .I(net_72624),
    .O(net_72624_cascademuxed)
  );
  CascadeMux t104 (
    .I(net_12612),
    .O(net_12612_cascademuxed)
  );
  CascadeMux t1040 (
    .I(net_72630),
    .O(net_72630_cascademuxed)
  );
  CascadeMux t1041 (
    .I(net_72642),
    .O(net_72642_cascademuxed)
  );
  CascadeMux t1042 (
    .I(net_72747),
    .O(net_72747_cascademuxed)
  );
  CascadeMux t1043 (
    .I(net_72753),
    .O(net_72753_cascademuxed)
  );
  CascadeMux t1044 (
    .I(net_72759),
    .O(net_72759_cascademuxed)
  );
  CascadeMux t1045 (
    .I(net_72765),
    .O(net_72765_cascademuxed)
  );
  CascadeMux t1046 (
    .I(net_72771),
    .O(net_72771_cascademuxed)
  );
  CascadeMux t1047 (
    .I(net_72777),
    .O(net_72777_cascademuxed)
  );
  CascadeMux t1048 (
    .I(net_72783),
    .O(net_72783_cascademuxed)
  );
  CascadeMux t1049 (
    .I(net_72789),
    .O(net_72789_cascademuxed)
  );
  CascadeMux t105 (
    .I(net_12618),
    .O(net_12618_cascademuxed)
  );
  CascadeMux t1050 (
    .I(net_72870),
    .O(net_72870_cascademuxed)
  );
  CascadeMux t1051 (
    .I(net_72993),
    .O(net_72993_cascademuxed)
  );
  CascadeMux t1052 (
    .I(net_73029),
    .O(net_73029_cascademuxed)
  );
  CascadeMux t1053 (
    .I(net_73116),
    .O(net_73116_cascademuxed)
  );
  CascadeMux t1054 (
    .I(net_73122),
    .O(net_73122_cascademuxed)
  );
  CascadeMux t1055 (
    .I(net_73128),
    .O(net_73128_cascademuxed)
  );
  CascadeMux t1056 (
    .I(net_73134),
    .O(net_73134_cascademuxed)
  );
  CascadeMux t1057 (
    .I(net_73140),
    .O(net_73140_cascademuxed)
  );
  CascadeMux t1058 (
    .I(net_73146),
    .O(net_73146_cascademuxed)
  );
  CascadeMux t1059 (
    .I(net_73275),
    .O(net_73275_cascademuxed)
  );
  CascadeMux t1060 (
    .I(net_73386),
    .O(net_73386_cascademuxed)
  );
  CascadeMux t1061 (
    .I(net_73404),
    .O(net_73404_cascademuxed)
  );
  CascadeMux t1062 (
    .I(net_73497),
    .O(net_73497_cascademuxed)
  );
  CascadeMux t1063 (
    .I(net_73521),
    .O(net_73521_cascademuxed)
  );
  CascadeMux t1064 (
    .I(net_73608),
    .O(net_73608_cascademuxed)
  );
  CascadeMux t1065 (
    .I(net_73626),
    .O(net_73626_cascademuxed)
  );
  CascadeMux t1066 (
    .I(net_73731),
    .O(net_73731_cascademuxed)
  );
  CascadeMux t1067 (
    .I(net_73737),
    .O(net_73737_cascademuxed)
  );
  CascadeMux t1068 (
    .I(net_73743),
    .O(net_73743_cascademuxed)
  );
  CascadeMux t1069 (
    .I(net_73749),
    .O(net_73749_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t107 (
    .carryinitin(),
    .carryinitout(t106)
  );
  CascadeMux t1070 (
    .I(net_73755),
    .O(net_73755_cascademuxed)
  );
  CascadeMux t1071 (
    .I(net_73761),
    .O(net_73761_cascademuxed)
  );
  CascadeMux t1072 (
    .I(net_73767),
    .O(net_73767_cascademuxed)
  );
  CascadeMux t1073 (
    .I(net_73773),
    .O(net_73773_cascademuxed)
  );
  CascadeMux t1074 (
    .I(net_73854),
    .O(net_73854_cascademuxed)
  );
  CascadeMux t1075 (
    .I(net_73878),
    .O(net_73878_cascademuxed)
  );
  CascadeMux t1076 (
    .I(net_79175),
    .O(net_79175_cascademuxed)
  );
  CascadeMux t1077 (
    .I(net_79415),
    .O(net_79415_cascademuxed)
  );
  CascadeMux t1078 (
    .I(net_79538),
    .O(net_79538_cascademuxed)
  );
  CascadeMux t1079 (
    .I(net_79655),
    .O(net_79655_cascademuxed)
  );
  CascadeMux t108 (
    .I(net_12699),
    .O(net_12699_cascademuxed)
  );
  CascadeMux t1080 (
    .I(net_79679),
    .O(net_79679_cascademuxed)
  );
  CascadeMux t1081 (
    .I(net_79685),
    .O(net_79685_cascademuxed)
  );
  CascadeMux t1082 (
    .I(net_79808),
    .O(net_79808_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t1084 (
    .carryinitin(),
    .carryinitout(t1083)
  );
  CascadeMux t1085 (
    .I(net_79937),
    .O(net_79937_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t1086 (
    .carryinitin(net_83771),
    .carryinitout(net_83815)
  );
  CascadeMux t1087 (
    .I(net_80048),
    .O(net_80048_cascademuxed)
  );
  CascadeMux t1088 (
    .I(net_80066),
    .O(net_80066_cascademuxed)
  );
  CascadeMux t1089 (
    .I(net_80177),
    .O(net_80177_cascademuxed)
  );
  CascadeMux t109 (
    .I(net_12705),
    .O(net_12705_cascademuxed)
  );
  CascadeMux t1090 (
    .I(net_80405),
    .O(net_80405_cascademuxed)
  );
  CascadeMux t1091 (
    .I(net_83252),
    .O(net_83252_cascademuxed)
  );
  CascadeMux t1092 (
    .I(net_83270),
    .O(net_83270_cascademuxed)
  );
  CascadeMux t1093 (
    .I(net_83399),
    .O(net_83399_cascademuxed)
  );
  CascadeMux t1094 (
    .I(net_83522),
    .O(net_83522_cascademuxed)
  );
  CascadeMux t1095 (
    .I(net_83627),
    .O(net_83627_cascademuxed)
  );
  CascadeMux t1096 (
    .I(net_83732),
    .O(net_83732_cascademuxed)
  );
  CascadeMux t1097 (
    .I(net_83738),
    .O(net_83738_cascademuxed)
  );
  CascadeMux t1098 (
    .I(net_83744),
    .O(net_83744_cascademuxed)
  );
  CascadeMux t1099 (
    .I(net_83750),
    .O(net_83750_cascademuxed)
  );
  CascadeMux t11 (
    .I(net_6967),
    .O(net_6967_cascademuxed)
  );
  CascadeMux t110 (
    .I(net_12711),
    .O(net_12711_cascademuxed)
  );
  CascadeMux t1100 (
    .I(net_83756),
    .O(net_83756_cascademuxed)
  );
  CascadeMux t1101 (
    .I(net_83762),
    .O(net_83762_cascademuxed)
  );
  CascadeMux t1102 (
    .I(net_83768),
    .O(net_83768_cascademuxed)
  );
  CascadeMux t1103 (
    .I(net_83774),
    .O(net_83774_cascademuxed)
  );
  CascadeMux t1104 (
    .I(net_83855),
    .O(net_83855_cascademuxed)
  );
  CascadeMux t1105 (
    .I(net_83861),
    .O(net_83861_cascademuxed)
  );
  CascadeMux t1106 (
    .I(net_83867),
    .O(net_83867_cascademuxed)
  );
  CascadeMux t1107 (
    .I(net_83897),
    .O(net_83897_cascademuxed)
  );
  CascadeMux t1108 (
    .I(net_83990),
    .O(net_83990_cascademuxed)
  );
  CascadeMux t1109 (
    .I(net_86948),
    .O(net_86948_cascademuxed)
  );
  CascadeMux t111 (
    .I(net_12717),
    .O(net_12717_cascademuxed)
  );
  CascadeMux t1110 (
    .I(net_86960),
    .O(net_86960_cascademuxed)
  );
  CascadeMux t1111 (
    .I(net_86972),
    .O(net_86972_cascademuxed)
  );
  CascadeMux t1112 (
    .I(net_87083),
    .O(net_87083_cascademuxed)
  );
  CascadeMux t1113 (
    .I(net_87113),
    .O(net_87113_cascademuxed)
  );
  CascadeMux t1114 (
    .I(net_87218),
    .O(net_87218_cascademuxed)
  );
  CascadeMux t1115 (
    .I(net_87236),
    .O(net_87236_cascademuxed)
  );
  CascadeMux t1116 (
    .I(net_87563),
    .O(net_87563_cascademuxed)
  );
  CascadeMux t1117 (
    .I(net_87575),
    .O(net_87575_cascademuxed)
  );
  CascadeMux t1118 (
    .I(net_91031),
    .O(net_91031_cascademuxed)
  );
  CascadeMux t1119 (
    .I(net_91067),
    .O(net_91067_cascademuxed)
  );
  CascadeMux t112 (
    .I(net_12723),
    .O(net_12723_cascademuxed)
  );
  LocalMux t1120 (
    .I(seg_4_11_sp4_v_b_25_16355),
    .O(seg_4_11_local_g2_1_20220)
  );
  Span4Mux_v2 t1121 (
    .I(seg_4_9_sp4_v_b_5_15867),
    .O(seg_4_11_sp4_v_b_25_16355)
  );
  Span4Mux_v4 t1122 (
    .I(seg_4_5_sp4_h_l_37_1178),
    .O(seg_4_9_sp4_v_b_5_15867)
  );
  LocalMux t1123 (
    .I(seg_8_5_sp4_h_r_18_30430),
    .O(seg_8_5_local_g0_2_34160)
  );
  Span4Mux_h1 t1124 (
    .I(seg_7_5_sp4_h_l_46_15731),
    .O(seg_8_5_sp4_h_r_18_30430)
  );
  Span4Mux_h4 t1125 (
    .I(seg_3_5_sp4_h_l_38_1184),
    .O(seg_7_5_sp4_h_l_46_15731)
  );
  LocalMux t1126 (
    .I(seg_1_13_sp4_r_v_b_8_8217),
    .O(seg_1_13_local_g2_0_8535)
  );
  Span4Mux_v4 t1127 (
    .I(seg_2_9_sp4_v_b_5_7624),
    .O(seg_1_13_sp4_r_v_b_8_8217)
  );
  Span4Mux_v4 t1128 (
    .I(seg_2_5_sp4_h_l_37_1195),
    .O(seg_2_9_sp4_v_b_5_7624)
  );
  LocalMux t1129 (
    .I(seg_1_13_sp4_r_v_b_4_8213),
    .O(seg_1_13_local_g1_4_8531)
  );
  CascadeMux t113 (
    .I(net_12729),
    .O(net_12729_cascademuxed)
  );
  Span4Mux_v4 t1130 (
    .I(seg_2_9_sp4_v_b_4_7625),
    .O(seg_1_13_sp4_r_v_b_4_8213)
  );
  Span4Mux_v4 t1131 (
    .I(seg_2_5_sp4_h_l_41_1199),
    .O(seg_2_9_sp4_v_b_4_7625)
  );
  LocalMux t1132 (
    .I(seg_2_13_sp4_v_b_11_8218),
    .O(seg_2_13_local_g1_3_12798)
  );
  Span4Mux_v4 t1133 (
    .I(seg_2_9_sp4_v_b_3_7622),
    .O(seg_2_13_sp4_v_b_11_8218)
  );
  Span4Mux_v4 t1134 (
    .I(seg_2_5_sp4_h_l_47_1206),
    .O(seg_2_9_sp4_v_b_3_7622)
  );
  LocalMux t1135 (
    .I(seg_1_13_sp4_v_b_11_2296),
    .O(seg_1_13_local_g0_3_8522)
  );
  Span4Mux_v4 t1136 (
    .I(seg_1_9_sp4_v_b_8_1441),
    .O(seg_1_13_sp4_v_b_11_2296)
  );
  Span4Mux_v4 t1137 (
    .I(seg_1_5_sp4_h_l_38_1210),
    .O(seg_1_9_sp4_v_b_8_1441)
  );
  LocalMux t1138 (
    .I(seg_1_13_sp4_v_b_22_2502),
    .O(seg_1_13_local_g0_6_8525)
  );
  Span4Mux_v3 t1139 (
    .I(seg_1_10_sp4_v_b_11_1650),
    .O(seg_1_13_sp4_v_b_22_2502)
  );
  CascadeMux t114 (
    .I(net_12735),
    .O(net_12735_cascademuxed)
  );
  Span4Mux_v4 t1140 (
    .I(seg_1_6_sp4_v_b_8_798),
    .O(seg_1_10_sp4_v_b_11_1650)
  );
  LocalMux t1141 (
    .I(seg_4_11_sp4_v_b_2_16112),
    .O(seg_4_11_local_g1_2_20213)
  );
  Span4Mux_v4 t1142 (
    .I(seg_4_7_sp4_h_l_39_1604),
    .O(seg_4_11_sp4_v_b_2_16112)
  );
  Span4Mux_h4 t1143 (
    .I(seg_0_7_sp4_v_b_2_804),
    .O(seg_4_7_sp4_h_l_39_1604)
  );
  LocalMux t1144 (
    .I(seg_7_10_sp4_r_v_b_8_30688),
    .O(seg_7_10_local_g2_0_30958)
  );
  Span4Mux_v4 t1145 (
    .I(seg_8_6_sp4_h_l_45_19692),
    .O(seg_7_10_sp4_r_v_b_8_30688)
  );
  Span4Mux_h4 t1146 (
    .I(seg_4_6_sp4_h_l_37_1384),
    .O(seg_8_6_sp4_h_l_45_19692)
  );
  LocalMux t1147 (
    .I(seg_7_13_sp4_r_v_b_21_31180),
    .O(seg_7_13_local_g3_5_31340)
  );
  Span4Mux_v3 t1148 (
    .I(seg_8_10_sp4_v_b_5_30683),
    .O(seg_7_13_sp4_r_v_b_21_31180)
  );
  Span4Mux_v4 t1149 (
    .I(seg_8_6_sp4_h_l_37_19682),
    .O(seg_8_10_sp4_v_b_5_30683)
  );
  CascadeMux t115 (
    .I(net_12741),
    .O(net_12741_cascademuxed)
  );
  Span4Mux_h4 t1150 (
    .I(seg_4_6_sp4_h_l_41_1418),
    .O(seg_8_6_sp4_h_l_37_19682)
  );
  LocalMux t1151 (
    .I(seg_8_5_sp4_r_v_b_13_34019),
    .O(seg_8_5_local_g2_5_34179)
  );
  Span4Mux_v1 t1152 (
    .I(seg_9_6_sp4_h_l_37_23513),
    .O(seg_8_5_sp4_r_v_b_13_34019)
  );
  Span4Mux_h4 t1153 (
    .I(seg_5_6_sp4_h_l_37_7608),
    .O(seg_9_6_sp4_h_l_37_23513)
  );
  Span4Mux_h4 t1154 (
    .I(seg_1_6_sp4_h_l_44_1423),
    .O(seg_5_6_sp4_h_l_37_7608)
  );
  LocalMux t1155 (
    .I(seg_2_6_sp4_h_r_32_1430),
    .O(seg_2_6_local_g3_0_11950)
  );
  LocalMux t1156 (
    .I(seg_7_7_sp4_h_r_28_23642),
    .O(seg_7_7_local_g3_4_30601)
  );
  Span4Mux_h2 t1157 (
    .I(seg_5_7_sp4_h_l_45_7765),
    .O(seg_7_7_sp4_h_r_28_23642)
  );
  Span4Mux_h4 t1158 (
    .I(seg_1_7_sp4_v_b_2_1019),
    .O(seg_5_7_sp4_h_l_45_7765)
  );
  LocalMux t1159 (
    .I(seg_5_11_sp4_v_b_0_19941),
    .O(seg_5_11_local_g1_0_24042)
  );
  Span4Mux_v4 t1160 (
    .I(seg_5_7_sp4_h_l_37_7755),
    .O(seg_5_11_sp4_v_b_0_19941)
  );
  Span4Mux_h4 t1161 (
    .I(seg_1_7_sp4_v_b_6_1023),
    .O(seg_5_7_sp4_h_l_37_7755)
  );
  LocalMux t1162 (
    .I(seg_7_8_sp4_h_r_24_23759),
    .O(seg_7_8_local_g3_0_30720)
  );
  Span4Mux_h2 t1163 (
    .I(seg_5_8_sp4_h_l_44_7913),
    .O(seg_7_8_sp4_h_r_24_23759)
  );
  Span4Mux_h4 t1164 (
    .I(seg_1_8_sp4_v_b_3_1228),
    .O(seg_5_8_sp4_h_l_44_7913)
  );
  LocalMux t1165 (
    .I(seg_7_11_sp4_r_v_b_11_30812),
    .O(seg_7_11_local_g2_3_31084)
  );
  Span4Mux_v4 t1166 (
    .I(seg_8_7_sp4_h_l_46_19808),
    .O(seg_7_11_sp4_r_v_b_11_30812)
  );
  Span4Mux_h4 t1167 (
    .I(seg_4_7_sp4_h_l_46_1595),
    .O(seg_8_7_sp4_h_l_46_19808)
  );
  Span4Mux_h4 t1168 (
    .I(seg_0_7_sp4_v_b_11_811),
    .O(seg_4_7_sp4_h_l_46_1595)
  );
  LocalMux t1169 (
    .I(seg_4_4_sp4_v_b_47_15628),
    .O(seg_4_4_local_g2_7_19365)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t117 (
    .carryinitin(),
    .carryinitout(t116)
  );
  Span4Mux_v3 t1170 (
    .I(seg_4_7_sp4_h_l_47_1594),
    .O(seg_4_4_sp4_v_b_47_15628)
  );
  LocalMux t1171 (
    .I(seg_3_5_sp4_v_b_33_11794),
    .O(seg_3_5_local_g2_1_15651)
  );
  Span4Mux_v2 t1172 (
    .I(seg_3_7_sp4_h_l_38_1598),
    .O(seg_3_5_sp4_v_b_33_11794)
  );
  LocalMux t1173 (
    .I(seg_2_6_sp4_v_b_15_7329),
    .O(seg_2_6_local_g1_7_11941)
  );
  Span4Mux_v1 t1174 (
    .I(seg_2_7_sp4_h_l_45_1618),
    .O(seg_2_6_sp4_v_b_15_7329)
  );
  LocalMux t1175 (
    .I(seg_7_7_sp4_h_r_39_19809),
    .O(seg_7_7_local_g3_7_30604)
  );
  Span4Mux_h3 t1176 (
    .I(seg_4_7_sp4_h_l_43_1636),
    .O(seg_7_7_sp4_h_r_39_19809)
  );
  LocalMux t1177 (
    .I(seg_8_4_sp4_h_r_37_23267),
    .O(seg_8_4_local_g3_5_34064)
  );
  Span4Mux_h3 t1178 (
    .I(seg_5_4_sp4_h_l_37_7314),
    .O(seg_8_4_sp4_h_r_37_23267)
  );
  Span4Mux_h4 t1179 (
    .I(seg_1_4_sp4_v_t_37_1227),
    .O(seg_5_4_sp4_h_l_37_7314)
  );
  CascadeMux t118 (
    .I(net_12822),
    .O(net_12822_cascademuxed)
  );
  LocalMux t1180 (
    .I(seg_5_8_sp4_h_r_9_23770),
    .O(seg_5_8_local_g1_1_23674)
  );
  Span4Mux_h0 t1181 (
    .I(seg_5_8_sp4_h_l_43_7910),
    .O(seg_5_8_sp4_h_r_9_23770)
  );
  Span4Mux_h4 t1182 (
    .I(seg_1_8_sp4_v_b_6_1233),
    .O(seg_5_8_sp4_h_l_43_7910)
  );
  LocalMux t1183 (
    .I(seg_5_8_sp4_h_r_5_23766),
    .O(seg_5_8_local_g0_5_23670)
  );
  Span4Mux_h0 t1184 (
    .I(seg_5_8_sp4_h_l_39_7906),
    .O(seg_5_8_sp4_h_r_5_23766)
  );
  Span4Mux_h4 t1185 (
    .I(seg_1_8_sp4_v_b_8_1235),
    .O(seg_5_8_sp4_h_l_39_7906)
  );
  LocalMux t1186 (
    .I(seg_5_8_sp4_v_b_33_19825),
    .O(seg_5_8_local_g2_1_23682)
  );
  Span4Mux_v2 t1187 (
    .I(seg_5_6_sp4_h_l_41_7614),
    .O(seg_5_8_sp4_v_b_33_19825)
  );
  Span4Mux_h4 t1188 (
    .I(seg_1_6_sp4_v_t_41_1645),
    .O(seg_5_6_sp4_h_l_41_7614)
  );
  LocalMux t1189 (
    .I(seg_4_5_sp4_v_b_37_15741),
    .O(seg_4_5_local_g3_5_19494)
  );
  CascadeMux t119 (
    .I(net_12828),
    .O(net_12828_cascademuxed)
  );
  Span4Mux_v3 t1190 (
    .I(seg_4_8_sp4_h_l_37_1801),
    .O(seg_4_5_sp4_v_b_37_15741)
  );
  LocalMux t1191 (
    .I(seg_7_2_sp4_v_b_25_26713),
    .O(seg_7_2_local_g3_1_29983)
  );
  Span4Mux_v2 t1192 (
    .I(seg_7_4_sp4_v_t_36_27127),
    .O(seg_7_2_sp4_v_b_25_26713)
  );
  Span4Mux_v4 t1193 (
    .I(seg_7_8_sp4_h_l_36_16098),
    .O(seg_7_4_sp4_v_t_36_27127)
  );
  Span4Mux_h4 t1194 (
    .I(seg_3_8_sp4_h_l_36_1805),
    .O(seg_7_8_sp4_h_l_36_16098)
  );
  LocalMux t1195 (
    .I(seg_10_5_sp4_r_v_b_38_41928),
    .O(seg_10_5_local_g2_6_41842)
  );
  Span4Mux_v3 t1196 (
    .I(seg_11_8_sp4_h_l_38_30795),
    .O(seg_10_5_sp4_r_v_b_38_41928)
  );
  Span4Mux_h4 t1197 (
    .I(seg_7_8_sp4_h_l_37_16097),
    .O(seg_11_8_sp4_h_l_38_30795)
  );
  Span4Mux_h4 t1198 (
    .I(seg_3_8_sp4_h_l_44_1814),
    .O(seg_7_8_sp4_h_l_37_16097)
  );
  LocalMux t1199 (
    .I(seg_1_5_sp4_v_b_42_1232),
    .O(seg_1_5_local_g2_2_7361)
  );
  CascadeMux t12 (
    .I(net_6979),
    .O(net_6979_cascademuxed)
  );
  CascadeMux t120 (
    .I(net_12840),
    .O(net_12840_cascademuxed)
  );
  LocalMux t1200 (
    .I(seg_8_2_sp4_v_b_29_29940),
    .O(seg_8_2_local_g3_5_33818)
  );
  Span4Mux_v2 t1201 (
    .I(seg_8_4_sp4_h_l_40_19443),
    .O(seg_8_2_sp4_v_b_29_29940)
  );
  Span4Mux_h4 t1202 (
    .I(seg_4_4_sp4_h_l_39_980),
    .O(seg_8_4_sp4_h_l_40_19443)
  );
  Span4Mux_h4 t1203 (
    .I(seg_0_4_sp4_v_t_39_1031),
    .O(seg_4_4_sp4_h_l_39_980)
  );
  LocalMux t1204 (
    .I(seg_3_5_sp4_r_v_b_18_15500),
    .O(seg_3_5_local_g3_2_15660)
  );
  Span4Mux_v1 t1205 (
    .I(seg_4_6_sp4_h_l_42_1429),
    .O(seg_3_5_sp4_r_v_b_18_15500)
  );
  Span4Mux_h4 t1206 (
    .I(seg_0_6_sp4_v_t_39_1447),
    .O(seg_4_6_sp4_h_l_42_1429)
  );
  LocalMux t1207 (
    .I(seg_7_1_sp4_r_v_b_44_29944),
    .O(seg_7_1_local_g3_4_29823)
  );
  Span4Mux_v3 t1208 (
    .I(seg_8_4_sp4_h_l_44_19447),
    .O(seg_7_1_sp4_r_v_b_44_29944)
  );
  Span4Mux_h4 t1209 (
    .I(seg_4_4_sp4_h_l_36_969),
    .O(seg_8_4_sp4_h_l_44_19447)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t121 (
    .carryinitin(net_16692),
    .carryinitout(net_16736)
  );
  Span4Mux_h4 t1210 (
    .I(seg_0_4_sp4_v_t_45_1037),
    .O(seg_4_4_sp4_h_l_36_969)
  );
  LocalMux t1211 (
    .I(seg_1_13_sp4_v_b_16_2496),
    .O(seg_1_13_local_g0_0_8519)
  );
  Span4Mux_v3 t1212 (
    .I(seg_1_10_sp4_h_l_40_2273),
    .O(seg_1_13_sp4_v_b_16_2496)
  );
  LocalMux t1213 (
    .I(seg_2_13_sp4_h_r_19_8645),
    .O(seg_2_13_local_g0_3_12790)
  );
  Span4Mux_h1 t1214 (
    .I(seg_1_13_sp4_v_b_0_2287),
    .O(seg_2_13_sp4_h_r_19_8645)
  );
  LocalMux t1215 (
    .I(seg_1_13_sp4_v_b_2_2289),
    .O(seg_1_13_local_g1_2_8529)
  );
  LocalMux t1216 (
    .I(seg_1_13_sp4_v_b_6_2293),
    .O(seg_1_13_local_g1_6_8533)
  );
  LocalMux t1217 (
    .I(seg_1_13_sp4_v_b_8_2295),
    .O(seg_1_13_local_g1_0_8527)
  );
  LocalMux t1218 (
    .I(seg_8_13_sp4_h_r_43_24382),
    .O(seg_8_13_local_g2_3_35161)
  );
  Span4Mux_h3 t1219 (
    .I(seg_5_13_sp4_h_l_47_8639),
    .O(seg_8_13_sp4_h_r_43_24382)
  );
  CascadeMux t122 (
    .I(net_12945),
    .O(net_12945_cascademuxed)
  );
  Span4Mux_h4 t1220 (
    .I(seg_1_13_sp4_v_b_10_2297),
    .O(seg_5_13_sp4_h_l_47_8639)
  );
  LocalMux t1221 (
    .I(seg_4_11_sp4_h_r_2_20301),
    .O(seg_4_11_local_g0_2_20205)
  );
  Span4Mux_h0 t1222 (
    .I(seg_4_11_sp4_h_l_46_2447),
    .O(seg_4_11_sp4_h_r_2_20301)
  );
  Span4Mux_h4 t1223 (
    .I(seg_0_11_sp4_v_b_5_1656),
    .O(seg_4_11_sp4_h_l_46_2447)
  );
  LocalMux t1224 (
    .I(seg_4_11_sp4_h_r_1_20298),
    .O(seg_4_11_local_g0_1_20204)
  );
  Span4Mux_h0 t1225 (
    .I(seg_4_11_sp4_h_l_36_2445),
    .O(seg_4_11_sp4_h_r_1_20298)
  );
  Span4Mux_h4 t1226 (
    .I(seg_0_11_sp4_v_b_7_1658),
    .O(seg_4_11_sp4_h_l_36_2445)
  );
  LocalMux t1227 (
    .I(seg_8_11_sp4_h_r_4_34996),
    .O(seg_8_11_local_g1_4_34908)
  );
  Span4Mux_h0 t1228 (
    .I(seg_8_11_sp4_h_l_45_20307),
    .O(seg_8_11_sp4_h_r_4_34996)
  );
  Span4Mux_h4 t1229 (
    .I(seg_4_11_sp4_h_l_37_2444),
    .O(seg_8_11_sp4_h_l_45_20307)
  );
  CascadeMux t123 (
    .I(net_12951),
    .O(net_12951_cascademuxed)
  );
  LocalMux t1230 (
    .I(seg_7_10_sp4_r_v_b_19_30809),
    .O(seg_7_10_local_g3_3_30969)
  );
  Span4Mux_v1 t1231 (
    .I(seg_8_11_sp4_h_l_43_20305),
    .O(seg_7_10_sp4_r_v_b_19_30809)
  );
  Span4Mux_h4 t1232 (
    .I(seg_4_11_sp4_h_l_47_2446),
    .O(seg_8_11_sp4_h_l_43_20305)
  );
  LocalMux t1233 (
    .I(seg_7_10_sp4_v_b_12_27433),
    .O(seg_7_10_local_g0_4_30946)
  );
  Span4Mux_v1 t1234 (
    .I(seg_7_11_sp4_h_l_36_16467),
    .O(seg_7_10_sp4_v_b_12_27433)
  );
  Span4Mux_h4 t1235 (
    .I(seg_3_11_sp4_h_l_36_2448),
    .O(seg_7_11_sp4_h_l_36_16467)
  );
  LocalMux t1236 (
    .I(seg_5_11_sp4_h_r_23_20299),
    .O(seg_5_11_local_g1_7_24049)
  );
  Span4Mux_h1 t1237 (
    .I(seg_4_11_sp4_h_l_39_2456),
    .O(seg_5_11_sp4_h_r_23_20299)
  );
  LocalMux t1238 (
    .I(seg_7_11_sp4_h_r_37_20297),
    .O(seg_7_11_local_g2_5_31086)
  );
  Span4Mux_h3 t1239 (
    .I(seg_4_11_sp4_h_l_41_2478),
    .O(seg_7_11_sp4_h_r_37_20297)
  );
  CascadeMux t124 (
    .I(net_12957),
    .O(net_12957_cascademuxed)
  );
  LocalMux t1240 (
    .I(seg_9_10_sp4_v_b_16_34637),
    .O(seg_9_10_local_g0_0_38604)
  );
  Span4Mux_v1 t1241 (
    .I(seg_9_11_sp4_h_l_40_24135),
    .O(seg_9_10_sp4_v_b_16_34637)
  );
  Span4Mux_h4 t1242 (
    .I(seg_5_11_sp4_h_l_39_8347),
    .O(seg_9_11_sp4_h_l_40_24135)
  );
  Span4Mux_h4 t1243 (
    .I(seg_1_11_sp4_h_l_46_2485),
    .O(seg_5_11_sp4_h_l_39_8347)
  );
  LocalMux t1244 (
    .I(seg_8_13_sp4_v_b_26_31297),
    .O(seg_8_13_local_g3_2_35168)
  );
  Span4Mux_v2 t1245 (
    .I(seg_8_11_sp4_h_l_44_20308),
    .O(seg_8_13_sp4_v_b_26_31297)
  );
  Span4Mux_h4 t1246 (
    .I(seg_4_11_sp4_h_l_43_2488),
    .O(seg_8_11_sp4_h_l_44_20308)
  );
  LocalMux t1247 (
    .I(seg_7_11_sp4_h_r_46_20300),
    .O(seg_7_11_local_g2_6_31087)
  );
  Span4Mux_h3 t1248 (
    .I(seg_4_11_sp4_h_l_45_2490),
    .O(seg_7_11_sp4_h_r_46_20300)
  );
  LocalMux t1249 (
    .I(seg_7_10_sp4_v_b_29_27539),
    .O(seg_7_10_local_g2_5_30963)
  );
  CascadeMux t125 (
    .I(net_12975),
    .O(net_12975_cascademuxed)
  );
  Span4Mux_v2 t1250 (
    .I(seg_7_12_sp4_h_l_40_16596),
    .O(seg_7_10_sp4_v_b_29_27539)
  );
  Span4Mux_h4 t1251 (
    .I(seg_3_12_sp4_h_l_40_2660),
    .O(seg_7_12_sp4_h_l_40_16596)
  );
  LocalMux t1252 (
    .I(seg_7_10_sp4_v_b_33_27543),
    .O(seg_7_10_local_g3_1_30967)
  );
  Span4Mux_v2 t1253 (
    .I(seg_7_12_sp4_h_l_44_16600),
    .O(seg_7_10_sp4_v_b_33_27543)
  );
  Span4Mux_h4 t1254 (
    .I(seg_3_12_sp4_h_l_44_2665),
    .O(seg_7_12_sp4_h_l_44_16600)
  );
  LocalMux t1255 (
    .I(seg_9_7_sp4_v_b_17_34269),
    .O(seg_9_7_local_g0_1_38236)
  );
  Span4Mux_v1 t1256 (
    .I(seg_9_8_sp4_h_l_41_23765),
    .O(seg_9_7_sp4_v_b_17_34269)
  );
  Span4Mux_h4 t1257 (
    .I(seg_5_8_sp4_h_l_41_7908),
    .O(seg_9_8_sp4_h_l_41_23765)
  );
  Span4Mux_h4 t1258 (
    .I(seg_1_8_sp4_v_t_46_2086),
    .O(seg_5_8_sp4_h_l_41_7908)
  );
  LocalMux t1259 (
    .I(seg_9_10_sp4_h_r_2_38702),
    .O(seg_9_10_local_g1_2_38614)
  );
  Span4Mux_h0 t1260 (
    .I(seg_9_10_sp4_h_l_43_24013),
    .O(seg_9_10_sp4_h_r_2_38702)
  );
  Span4Mux_h4 t1261 (
    .I(seg_5_10_sp4_h_l_43_8204),
    .O(seg_9_10_sp4_h_l_43_24013)
  );
  Span4Mux_h4 t1262 (
    .I(seg_1_10_sp4_v_t_36_2492),
    .O(seg_5_10_sp4_h_l_43_8204)
  );
  LocalMux t1263 (
    .I(seg_9_9_sp4_v_b_20_34518),
    .O(seg_9_9_local_g0_4_38485)
  );
  Span4Mux_v1 t1264 (
    .I(seg_9_10_sp4_h_l_38_24010),
    .O(seg_9_9_sp4_v_b_20_34518)
  );
  Span4Mux_h4 t1265 (
    .I(seg_5_10_sp4_h_l_37_8196),
    .O(seg_9_10_sp4_h_l_38_24010)
  );
  Span4Mux_h4 t1266 (
    .I(seg_1_10_sp4_v_t_42_2498),
    .O(seg_5_10_sp4_h_l_37_8196)
  );
  LocalMux t1267 (
    .I(seg_8_11_sp4_h_r_38_24133),
    .O(seg_8_11_local_g3_6_34926)
  );
  Span4Mux_h3 t1268 (
    .I(seg_5_11_sp4_h_l_42_8352),
    .O(seg_8_11_sp4_h_r_38_24133)
  );
  Span4Mux_h4 t1269 (
    .I(seg_1_11_sp4_v_t_39_2703),
    .O(seg_5_11_sp4_h_l_42_8352)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t127 (
    .carryinitin(),
    .carryinitout(t126)
  );
  LocalMux t1270 (
    .I(seg_8_2_sp4_v_b_39_30067),
    .O(seg_8_2_local_g2_7_33812)
  );
  Span4Mux_v3 t1271 (
    .I(seg_8_5_sp4_h_l_39_19563),
    .O(seg_8_2_sp4_v_b_39_30067)
  );
  Span4Mux_h4 t1272 (
    .I(seg_4_5_sp4_h_l_43_1222),
    .O(seg_8_5_sp4_h_l_39_19563)
  );
  Span4Mux_h4 t1273 (
    .I(seg_0_5_sp4_v_t_36_1238),
    .O(seg_4_5_sp4_h_l_43_1222)
  );
  Span4Mux_v4 t1274 (
    .I(seg_0_9_sp4_v_t_36_2088),
    .O(seg_0_5_sp4_v_t_36_1238)
  );
  LocalMux t1275 (
    .I(seg_9_10_sp4_h_r_19_34875),
    .O(seg_9_10_local_g1_3_38615)
  );
  Span4Mux_h1 t1276 (
    .I(seg_8_10_sp4_h_l_43_20182),
    .O(seg_9_10_sp4_h_r_19_34875)
  );
  Span4Mux_h4 t1277 (
    .I(seg_4_10_sp4_h_l_47_2240),
    .O(seg_8_10_sp4_h_l_43_20182)
  );
  Span4Mux_h4 t1278 (
    .I(seg_0_10_sp4_v_t_47_2309),
    .O(seg_4_10_sp4_h_l_47_2240)
  );
  LocalMux t1279 (
    .I(seg_9_9_sp4_h_r_22_34747),
    .O(seg_9_9_local_g0_6_38487)
  );
  CascadeMux t128 (
    .I(net_13068),
    .O(net_13068_cascademuxed)
  );
  Span4Mux_h1 t1280 (
    .I(seg_8_9_sp4_v_t_43_31055),
    .O(seg_9_9_sp4_h_r_22_34747)
  );
  Span4Mux_v4 t1281 (
    .I(seg_8_13_sp4_h_l_37_20543),
    .O(seg_8_9_sp4_v_t_43_31055)
  );
  Span4Mux_h4 t1282 (
    .I(seg_4_13_sp4_h_l_37_2861),
    .O(seg_8_13_sp4_h_l_37_20543)
  );
  LocalMux t1283 (
    .I(seg_4_5_sp4_h_r_31_11906),
    .O(seg_4_5_local_g3_7_19496)
  );
  Span4Mux_h2 t1284 (
    .I(seg_2_5_sp4_v_t_39_7623),
    .O(seg_4_5_sp4_h_r_31_11906)
  );
  Span4Mux_v4 t1285 (
    .I(seg_2_9_sp4_v_t_43_8215),
    .O(seg_2_5_sp4_v_t_39_7623)
  );
  Span4Mux_v4 t1286 (
    .I(seg_2_13_sp4_h_l_37_2878),
    .O(seg_2_9_sp4_v_t_43_8215)
  );
  LocalMux t1287 (
    .I(seg_5_8_sp4_v_b_22_19704),
    .O(seg_5_8_local_g0_6_23671)
  );
  Span4Mux_v1 t1288 (
    .I(seg_5_9_sp4_v_t_46_20196),
    .O(seg_5_8_sp4_v_b_22_19704)
  );
  Span4Mux_v4 t1289 (
    .I(seg_5_13_sp4_h_l_46_8640),
    .O(seg_5_9_sp4_v_t_46_20196)
  );
  CascadeMux t129 (
    .I(net_13074),
    .O(net_13074_cascademuxed)
  );
  Span4Mux_h4 t1290 (
    .I(seg_1_13_sp4_h_l_38_2893),
    .O(seg_5_13_sp4_h_l_46_8640)
  );
  LocalMux t1291 (
    .I(seg_10_10_sp4_h_r_18_38707),
    .O(seg_10_10_local_g0_2_42437)
  );
  Span4Mux_h1 t1292 (
    .I(seg_9_10_sp4_h_l_41_24011),
    .O(seg_10_10_sp4_h_r_18_38707)
  );
  Span4Mux_h4 t1293 (
    .I(seg_5_10_sp4_h_l_36_8197),
    .O(seg_9_10_sp4_h_l_41_24011)
  );
  Span4Mux_h4 t1294 (
    .I(seg_1_10_sp4_v_t_45_2501),
    .O(seg_5_10_sp4_h_l_36_8197)
  );
  LocalMux t1295 (
    .I(seg_1_8_sp4_v_b_46_1859),
    .O(seg_1_8_local_g2_6_7806)
  );
  Span4Mux_v3 t1296 (
    .I(seg_1_11_sp4_v_t_38_2702),
    .O(seg_1_8_sp4_v_b_46_1859)
  );
  LocalMux t1297 (
    .I(seg_1_5_sp4_h_r_3_7466),
    .O(seg_1_5_local_g0_3_7346)
  );
  Span4Mux_h0 t1298 (
    .I(seg_1_5_sp4_v_t_38_1434),
    .O(seg_1_5_sp4_h_r_3_7466)
  );
  Span4Mux_v4 t1299 (
    .I(seg_1_9_sp4_v_t_38_2288),
    .O(seg_1_5_sp4_v_t_38_1434)
  );
  CascadeMux t13 (
    .I(net_7084),
    .O(net_7084_cascademuxed)
  );
  CascadeMux t130 (
    .I(net_13080),
    .O(net_13080_cascademuxed)
  );
  LocalMux t1300 (
    .I(seg_3_10_sp4_h_r_43_2282),
    .O(seg_3_10_local_g3_3_16276)
  );
  Span4Mux_h3 t1301 (
    .I(seg_0_10_sp4_v_t_36_2298),
    .O(seg_3_10_sp4_h_r_43_2282)
  );
  LocalMux t1302 (
    .I(seg_4_17_sp4_v_b_34_17104),
    .O(seg_4_17_local_g3_2_20967)
  );
  Span4Mux_v2 t1303 (
    .I(seg_4_15_sp4_h_l_47_3300),
    .O(seg_4_17_sp4_v_b_34_17104)
  );
  LocalMux t1304 (
    .I(seg_2_14_sp4_r_v_b_14_12772),
    .O(seg_2_14_local_g2_6_12932)
  );
  Span4Mux_v1 t1305 (
    .I(seg_3_15_sp4_h_l_38_3304),
    .O(seg_2_14_sp4_r_v_b_14_12772)
  );
  LocalMux t1306 (
    .I(seg_7_16_sp4_v_b_47_28260),
    .O(seg_7_16_local_g3_7_31711)
  );
  Span4Mux_v1 t1307 (
    .I(seg_7_15_sp4_h_l_40_16965),
    .O(seg_7_16_sp4_v_b_47_28260)
  );
  Span4Mux_h4 t1308 (
    .I(seg_3_15_sp4_h_l_40_3306),
    .O(seg_7_15_sp4_h_l_40_16965)
  );
  LocalMux t1309 (
    .I(seg_7_16_sp4_v_b_37_28250),
    .O(seg_7_16_local_g3_5_31709)
  );
  CascadeMux t131 (
    .I(net_13086),
    .O(net_13086_cascademuxed)
  );
  Span4Mux_v1 t1310 (
    .I(seg_7_15_sp4_h_l_42_16967),
    .O(seg_7_16_sp4_v_b_37_28250)
  );
  Span4Mux_h4 t1311 (
    .I(seg_3_15_sp4_h_l_42_3308),
    .O(seg_7_15_sp4_h_l_42_16967)
  );
  LocalMux t1312 (
    .I(seg_4_17_sp4_v_b_25_17093),
    .O(seg_4_17_local_g2_1_20958)
  );
  Span4Mux_v2 t1313 (
    .I(seg_4_15_sp4_h_l_45_3344),
    .O(seg_4_17_sp4_v_b_25_17093)
  );
  LocalMux t1314 (
    .I(seg_7_16_sp4_h_r_24_24743),
    .O(seg_7_16_local_g2_0_31696)
  );
  Span4Mux_h2 t1315 (
    .I(seg_5_16_sp4_h_l_41_9084),
    .O(seg_7_16_sp4_h_r_24_24743)
  );
  Span4Mux_h4 t1316 (
    .I(seg_1_16_sp4_v_b_10_2920),
    .O(seg_5_16_sp4_h_l_41_9084)
  );
  LocalMux t1317 (
    .I(seg_7_16_sp4_h_r_37_20912),
    .O(seg_7_16_local_g2_5_31701)
  );
  Span4Mux_h3 t1318 (
    .I(seg_4_16_sp4_h_l_44_3551),
    .O(seg_7_16_sp4_h_r_37_20912)
  );
  Span4Mux_h4 t1319 (
    .I(seg_0_16_sp4_v_b_9_2720),
    .O(seg_4_16_sp4_h_l_44_3551)
  );
  CascadeMux t132 (
    .I(net_13203),
    .O(net_13203_cascademuxed)
  );
  LocalMux t1320 (
    .I(seg_4_17_sp4_h_r_6_21043),
    .O(seg_4_17_local_g1_6_20955)
  );
  Span4Mux_h0 t1321 (
    .I(seg_4_17_sp4_h_l_47_3714),
    .O(seg_4_17_sp4_h_r_6_21043)
  );
  Span4Mux_h4 t1322 (
    .I(seg_0_17_sp4_v_b_4_2926),
    .O(seg_4_17_sp4_h_l_47_3714)
  );
  LocalMux t1323 (
    .I(seg_3_14_sp4_v_b_25_12893),
    .O(seg_3_14_local_g2_1_16758)
  );
  Span4Mux_v2 t1324 (
    .I(seg_3_16_sp4_h_l_42_3514),
    .O(seg_3_14_sp4_v_b_25_12893)
  );
  LocalMux t1325 (
    .I(seg_1_15_sp4_v_b_24_3137),
    .O(seg_1_15_local_g2_0_8829)
  );
  LocalMux t1326 (
    .I(seg_1_12_sp4_v_b_16_2290),
    .O(seg_1_12_local_g1_0_8380)
  );
  Span4Mux_v1 t1327 (
    .I(seg_1_13_sp4_v_t_39_3139),
    .O(seg_1_12_sp4_v_b_16_2290)
  );
  LocalMux t1328 (
    .I(seg_1_9_sp4_v_b_45_2085),
    .O(seg_1_9_local_g3_5_7960)
  );
  Span4Mux_v3 t1329 (
    .I(seg_1_12_sp4_v_t_40_2913),
    .O(seg_1_9_sp4_v_b_45_2085)
  );
  CascadeMux t133 (
    .I(net_13227),
    .O(net_13227_cascademuxed)
  );
  LocalMux t1330 (
    .I(seg_2_14_sp4_h_r_26_3100),
    .O(seg_2_14_local_g2_2_12928)
  );
  Span4Mux_h2 t1331 (
    .I(seg_0_14_sp4_v_t_39_3151),
    .O(seg_2_14_sp4_h_r_26_3100)
  );
  LocalMux t1332 (
    .I(seg_2_14_sp4_h_r_25_3089),
    .O(seg_2_14_local_g2_1_12927)
  );
  Span4Mux_h2 t1333 (
    .I(seg_0_14_sp4_v_t_45_3157),
    .O(seg_2_14_sp4_h_r_25_3089)
  );
  LocalMux t1334 (
    .I(seg_1_12_sp4_h_r_19_2696),
    .O(seg_1_12_local_g1_3_8383)
  );
  Span4Mux_h1 t1335 (
    .I(seg_0_12_sp4_v_t_43_2719),
    .O(seg_1_12_sp4_h_r_19_2696)
  );
  LocalMux t1336 (
    .I(seg_1_12_sp4_h_r_12_2653),
    .O(seg_1_12_local_g1_4_8384)
  );
  Span4Mux_h1 t1337 (
    .I(seg_0_12_sp4_v_t_45_2721),
    .O(seg_1_12_sp4_h_r_12_2653)
  );
  LocalMux t1338 (
    .I(seg_2_14_sp4_v_b_45_8805),
    .O(seg_2_14_local_g2_5_12931)
  );
  Span4Mux_v3 t1339 (
    .I(seg_2_17_sp4_h_l_39_3731),
    .O(seg_2_14_sp4_v_b_45_8805)
  );
  CascadeMux t134 (
    .I(net_13233),
    .O(net_13233_cascademuxed)
  );
  LocalMux t1340 (
    .I(seg_4_15_sp4_v_b_34_16858),
    .O(seg_4_15_local_g2_2_20713)
  );
  Span4Mux_v2 t1341 (
    .I(seg_4_17_sp4_h_l_41_3746),
    .O(seg_4_15_sp4_v_b_34_16858)
  );
  LocalMux t1342 (
    .I(seg_4_14_sp4_v_b_45_16856),
    .O(seg_4_14_local_g3_5_20601)
  );
  Span4Mux_v3 t1343 (
    .I(seg_4_17_sp4_h_l_45_3758),
    .O(seg_4_14_sp4_v_b_45_16856)
  );
  LocalMux t1344 (
    .I(seg_1_15_sp4_v_b_41_3351),
    .O(seg_1_15_local_g2_1_8830)
  );
  LocalMux t1345 (
    .I(seg_5_15_sp4_h_r_1_24621),
    .O(seg_5_15_local_g1_1_24535)
  );
  Span4Mux_h0 t1346 (
    .I(seg_5_15_sp4_h_l_47_8933),
    .O(seg_5_15_sp4_h_r_1_24621)
  );
  Span4Mux_h4 t1347 (
    .I(seg_1_15_sp4_v_t_40_3556),
    .O(seg_5_15_sp4_h_l_47_8933)
  );
  LocalMux t1348 (
    .I(seg_5_15_sp4_h_r_4_24626),
    .O(seg_5_15_local_g1_4_24538)
  );
  Span4Mux_h0 t1349 (
    .I(seg_5_15_sp4_h_l_41_8937),
    .O(seg_5_15_sp4_h_r_4_24626)
  );
  CascadeMux t135 (
    .I(net_13356),
    .O(net_13356_cascademuxed)
  );
  Span4Mux_h4 t1350 (
    .I(seg_1_15_sp4_v_t_46_3562),
    .O(seg_5_15_sp4_h_l_41_8937)
  );
  LocalMux t1351 (
    .I(seg_1_14_sp4_h_r_22_3091),
    .O(seg_1_14_local_g1_6_8680)
  );
  Span4Mux_h1 t1352 (
    .I(seg_0_14_sp4_v_t_46_3158),
    .O(seg_1_14_sp4_h_r_22_3091)
  );
  LocalMux t1353 (
    .I(seg_2_15_sp4_h_r_30_3342),
    .O(seg_2_15_local_g2_6_13055)
  );
  Span4Mux_h2 t1354 (
    .I(seg_0_15_sp4_v_t_43_3365),
    .O(seg_2_15_sp4_h_r_30_3342)
  );
  LocalMux t1355 (
    .I(seg_4_16_sp4_v_b_24_16971),
    .O(seg_4_16_local_g2_0_20834)
  );
  Span4Mux_v2 t1356 (
    .I(seg_4_18_sp4_h_l_43_3965),
    .O(seg_4_16_sp4_v_b_24_16971)
  );
  LocalMux t1357 (
    .I(seg_1_15_sp4_v_b_46_3356),
    .O(seg_1_15_local_g2_6_8835)
  );
  LocalMux t1358 (
    .I(seg_1_16_sp4_v_b_37_3553),
    .O(seg_1_16_local_g3_5_8989)
  );
  LocalMux t1359 (
    .I(seg_1_15_sp4_h_r_11_8934),
    .O(seg_1_15_local_g1_3_8824)
  );
  CascadeMux t136 (
    .I(net_13479),
    .O(net_13479_cascademuxed)
  );
  Span4Mux_h0 t1360 (
    .I(seg_1_15_sp4_v_t_43_3559),
    .O(seg_1_15_sp4_h_r_11_8934)
  );
  LocalMux t1361 (
    .I(seg_1_16_sp4_v_b_29_3350),
    .O(seg_1_16_local_g2_5_8981)
  );
  LocalMux t1362 (
    .I(seg_1_16_sp4_v_b_33_3354),
    .O(seg_1_16_local_g2_1_8977)
  );
  LocalMux t1363 (
    .I(seg_2_15_sp4_h_r_29_3341),
    .O(seg_2_15_local_g3_5_13062)
  );
  Span4Mux_h2 t1364 (
    .I(seg_0_15_sp4_v_t_40_3362),
    .O(seg_2_15_sp4_h_r_29_3341)
  );
  LocalMux t1365 (
    .I(seg_7_18_sp4_r_v_b_22_31796),
    .O(seg_7_18_local_g3_6_31956)
  );
  Span4Mux_v1 t1366 (
    .I(seg_8_19_sp4_h_l_40_21288),
    .O(seg_7_18_sp4_r_v_b_22_31796)
  );
  Span4Mux_h4 t1367 (
    .I(seg_4_19_sp4_v_t_37_17586),
    .O(seg_8_19_sp4_h_l_40_21288)
  );
  Span4Mux_v4 t1368 (
    .I(seg_4_23_sp4_h_l_37_5039),
    .O(seg_4_19_sp4_v_t_37_17586)
  );
  LocalMux t1369 (
    .I(seg_7_19_sp4_h_r_24_25112),
    .O(seg_7_19_local_g2_0_32065)
  );
  CascadeMux t137 (
    .I(net_13560),
    .O(net_13560_cascademuxed)
  );
  Span4Mux_h2 t1370 (
    .I(seg_5_19_sp4_h_l_41_9525),
    .O(seg_7_19_sp4_h_r_24_25112)
  );
  Span4Mux_h4 t1371 (
    .I(seg_1_19_sp4_v_t_46_4433),
    .O(seg_5_19_sp4_h_l_41_9525)
  );
  LocalMux t1372 (
    .I(seg_1_17_sp4_v_b_47_3771),
    .O(seg_1_17_local_g2_7_9130)
  );
  Span4Mux_v3 t1373 (
    .I(seg_1_20_sp4_v_t_39_4653),
    .O(seg_1_17_sp4_v_b_47_3771)
  );
  LocalMux t1374 (
    .I(seg_5_19_sp4_h_r_6_25120),
    .O(seg_5_19_local_g0_6_25024)
  );
  Span4Mux_h0 t1375 (
    .I(seg_5_19_sp4_h_l_38_9524),
    .O(seg_5_19_sp4_h_r_6_25120)
  );
  Span4Mux_h4 t1376 (
    .I(seg_1_19_sp4_v_t_38_4425),
    .O(seg_5_19_sp4_h_l_38_9524)
  );
  LocalMux t1377 (
    .I(seg_7_19_sp4_h_r_29_25119),
    .O(seg_7_19_local_g2_5_32070)
  );
  Span4Mux_h2 t1378 (
    .I(seg_5_19_sp4_h_l_40_9526),
    .O(seg_7_19_sp4_h_r_29_25119)
  );
  Span4Mux_h4 t1379 (
    .I(seg_1_19_sp4_v_t_40_4427),
    .O(seg_5_19_sp4_h_l_40_9526)
  );
  CascadeMux t138 (
    .I(net_13596),
    .O(net_13596_cascademuxed)
  );
  LocalMux t1380 (
    .I(seg_4_19_sp4_h_r_42_9528),
    .O(seg_4_19_local_g2_2_21205)
  );
  Span4Mux_h3 t1381 (
    .I(seg_1_19_sp4_v_t_42_4429),
    .O(seg_4_19_sp4_h_r_42_9528)
  );
  LocalMux t1382 (
    .I(seg_7_19_sp4_h_r_33_25123),
    .O(seg_7_19_local_g3_1_32074)
  );
  Span4Mux_h2 t1383 (
    .I(seg_5_19_sp4_h_l_44_9530),
    .O(seg_7_19_sp4_h_r_33_25123)
  );
  Span4Mux_h4 t1384 (
    .I(seg_1_19_sp4_v_t_44_4431),
    .O(seg_5_19_sp4_h_l_44_9530)
  );
  LocalMux t1385 (
    .I(seg_7_19_sp4_r_v_b_15_31912),
    .O(seg_7_19_local_g2_7_32072)
  );
  Span4Mux_v1 t1386 (
    .I(seg_8_20_sp4_h_l_39_21408),
    .O(seg_7_19_sp4_r_v_b_15_31912)
  );
  Span4Mux_h4 t1387 (
    .I(seg_4_20_sp4_h_l_43_4419),
    .O(seg_8_20_sp4_h_l_39_21408)
  );
  Span4Mux_h4 t1388 (
    .I(seg_0_20_sp4_v_t_36_4435),
    .O(seg_4_20_sp4_h_l_43_4419)
  );
  LocalMux t1389 (
    .I(seg_2_18_sp4_r_v_b_35_13395),
    .O(seg_2_18_local_g2_3_13421)
  );
  CascadeMux t139 (
    .I(net_13959),
    .O(net_13959_cascademuxed)
  );
  Span4Mux_v2 t1390 (
    .I(seg_3_20_sp4_v_t_46_13887),
    .O(seg_2_18_sp4_r_v_b_35_13395)
  );
  Span4Mux_v4 t1391 (
    .I(seg_3_24_sp4_h_l_46_5260),
    .O(seg_3_20_sp4_v_t_46_13887)
  );
  LocalMux t1392 (
    .I(seg_1_14_sp4_v_b_31_2915),
    .O(seg_1_14_local_g2_7_8689)
  );
  Span4Mux_v2 t1393 (
    .I(seg_1_16_sp4_v_t_41_3765),
    .O(seg_1_14_sp4_v_b_31_2915)
  );
  Span4Mux_v4 t1394 (
    .I(seg_1_20_sp4_v_t_36_4650),
    .O(seg_1_16_sp4_v_t_41_3765)
  );
  LocalMux t1395 (
    .I(seg_1_14_sp4_v_b_26_2912),
    .O(seg_1_14_local_g2_2_8684)
  );
  Span4Mux_v2 t1396 (
    .I(seg_1_16_sp4_v_t_39_3763),
    .O(seg_1_14_sp4_v_b_26_2912)
  );
  Span4Mux_v4 t1397 (
    .I(seg_1_20_sp4_v_t_46_4660),
    .O(seg_1_16_sp4_v_t_39_3763)
  );
  LocalMux t1398 (
    .I(seg_3_21_sp4_h_r_26_9817),
    .O(seg_3_21_local_g2_2_17620)
  );
  Span4Mux_h2 t1399 (
    .I(seg_1_21_sp4_v_t_39_4880),
    .O(seg_3_21_sp4_h_r_26_9817)
  );
  CascadeMux t14 (
    .I(net_7090),
    .O(net_7090_cascademuxed)
  );
  CascadeMux t140 (
    .I(net_15137),
    .O(net_15137_cascademuxed)
  );
  LocalMux t1400 (
    .I(seg_1_18_sp4_h_r_10_9374),
    .O(seg_1_18_local_g0_2_9256)
  );
  Span4Mux_h0 t1401 (
    .I(seg_1_18_sp4_v_t_40_4200),
    .O(seg_1_18_sp4_h_r_10_9374)
  );
  Span4Mux_v4 t1402 (
    .I(seg_1_22_sp4_v_t_40_5091),
    .O(seg_1_18_sp4_v_t_40_4200)
  );
  LocalMux t1403 (
    .I(seg_2_18_sp4_h_r_22_9375),
    .O(seg_2_18_local_g0_6_13408)
  );
  Span4Mux_h1 t1404 (
    .I(seg_1_18_sp4_v_t_46_4206),
    .O(seg_2_18_sp4_h_r_22_9375)
  );
  Span4Mux_v4 t1405 (
    .I(seg_1_22_sp4_v_t_46_5097),
    .O(seg_1_18_sp4_v_t_46_4206)
  );
  LocalMux t1406 (
    .I(seg_1_14_sp4_v_b_33_2917),
    .O(seg_1_14_local_g2_1_8683)
  );
  Span4Mux_v2 t1407 (
    .I(seg_1_16_sp4_v_t_36_3760),
    .O(seg_1_14_sp4_v_b_33_2917)
  );
  Span4Mux_v4 t1408 (
    .I(seg_1_20_sp4_v_t_40_4654),
    .O(seg_1_16_sp4_v_t_36_3760)
  );
  LocalMux t1409 (
    .I(seg_3_20_sp4_h_r_33_9677),
    .O(seg_3_20_local_g3_1_17504)
  );
  CascadeMux t141 (
    .I(net_15143),
    .O(net_15143_cascademuxed)
  );
  Span4Mux_h2 t1410 (
    .I(seg_1_20_sp4_v_t_44_4658),
    .O(seg_3_20_sp4_h_r_33_9677)
  );
  LocalMux t1411 (
    .I(seg_4_20_sp4_v_b_21_17348),
    .O(seg_4_20_local_g0_5_21315)
  );
  Span4Mux_v1 t1412 (
    .I(seg_4_21_sp4_v_t_37_17832),
    .O(seg_4_20_sp4_v_b_21_17348)
  );
  Span4Mux_v4 t1413 (
    .I(seg_4_25_sp4_h_l_37_5453),
    .O(seg_4_21_sp4_v_t_37_17832)
  );
  LocalMux t1414 (
    .I(seg_2_20_sp4_v_b_23_9395),
    .O(seg_2_20_local_g0_7_13655)
  );
  Span4Mux_v1 t1415 (
    .I(seg_2_21_sp4_v_t_39_9975),
    .O(seg_2_20_sp4_v_b_23_9395)
  );
  Span4Mux_v4 t1416 (
    .I(seg_2_25_sp4_h_l_39_5472),
    .O(seg_2_21_sp4_v_t_39_9975)
  );
  LocalMux t1417 (
    .I(seg_4_20_sp4_v_b_15_17342),
    .O(seg_4_20_local_g0_7_21317)
  );
  Span4Mux_v1 t1418 (
    .I(seg_4_21_sp4_v_t_43_17838),
    .O(seg_4_20_sp4_v_b_15_17342)
  );
  Span4Mux_v4 t1419 (
    .I(seg_4_25_sp4_h_l_43_5497),
    .O(seg_4_21_sp4_v_t_43_17838)
  );
  CascadeMux t142 (
    .I(net_15149),
    .O(net_15149_cascademuxed)
  );
  LocalMux t1420 (
    .I(seg_4_22_sp4_v_b_39_17834),
    .O(seg_4_22_local_g2_7_21579)
  );
  Span4Mux_v3 t1421 (
    .I(seg_4_25_sp4_h_l_45_5499),
    .O(seg_4_22_sp4_v_b_39_17834)
  );
  LocalMux t1422 (
    .I(seg_1_20_sp4_v_b_24_4197),
    .O(seg_1_20_local_g2_0_9564)
  );
  Span4Mux_v2 t1423 (
    .I(seg_1_22_sp4_v_t_37_5088),
    .O(seg_1_20_sp4_v_b_24_4197)
  );
  LocalMux t1424 (
    .I(seg_1_20_sp4_v_b_22_3979),
    .O(seg_1_20_local_g0_6_9554)
  );
  Span4Mux_v1 t1425 (
    .I(seg_1_21_sp4_v_t_38_4879),
    .O(seg_1_20_sp4_v_b_22_3979)
  );
  LocalMux t1426 (
    .I(seg_1_21_sp4_v_b_34_4434),
    .O(seg_1_21_local_g3_2_9721)
  );
  Span4Mux_v2 t1427 (
    .I(seg_1_23_sp4_v_t_42_5299),
    .O(seg_1_21_sp4_v_b_34_4434)
  );
  LocalMux t1428 (
    .I(seg_1_20_sp4_v_b_12_3969),
    .O(seg_1_20_local_g1_4_9560)
  );
  Span4Mux_v1 t1429 (
    .I(seg_1_21_sp4_v_t_40_4881),
    .O(seg_1_20_sp4_v_b_12_3969)
  );
  CascadeMux t143 (
    .I(net_15155),
    .O(net_15155_cascademuxed)
  );
  LocalMux t1430 (
    .I(seg_2_22_sp4_h_r_3_13993),
    .O(seg_2_22_local_g0_3_13897)
  );
  Span4Mux_h0 t1431 (
    .I(seg_2_22_sp4_v_t_47_10130),
    .O(seg_2_22_sp4_h_r_3_13993)
  );
  Span4Mux_v4 t1432 (
    .I(seg_2_26_sp4_h_l_41_5683),
    .O(seg_2_22_sp4_v_t_47_10130)
  );
  LocalMux t1433 (
    .I(seg_2_23_sp4_h_r_17_10113),
    .O(seg_2_23_local_g1_1_14026)
  );
  Span4Mux_h1 t1434 (
    .I(seg_1_23_sp4_v_t_41_5298),
    .O(seg_2_23_sp4_h_r_17_10113)
  );
  LocalMux t1435 (
    .I(seg_2_19_sp4_h_r_12_9520),
    .O(seg_2_19_local_g0_4_13529)
  );
  Span4Mux_h1 t1436 (
    .I(seg_1_19_sp4_v_t_45_4432),
    .O(seg_2_19_sp4_h_r_12_9520)
  );
  Span4Mux_v4 t1437 (
    .I(seg_1_23_sp4_v_t_45_5302),
    .O(seg_1_19_sp4_v_t_45_4432)
  );
  LocalMux t1438 (
    .I(seg_2_20_sp4_h_r_13_9666),
    .O(seg_2_20_local_g0_5_13653)
  );
  Span4Mux_h1 t1439 (
    .I(seg_1_20_sp4_v_t_42_4656),
    .O(seg_2_20_sp4_h_r_13_9666)
  );
  CascadeMux t144 (
    .I(net_15173),
    .O(net_15173_cascademuxed)
  );
  Span4Mux_v4 t1440 (
    .I(seg_1_24_sp4_v_t_46_5511),
    .O(seg_1_20_sp4_v_t_42_4656)
  );
  LocalMux t1441 (
    .I(seg_1_23_sp4_v_b_42_5093),
    .O(seg_1_23_local_g3_2_10015)
  );
  LocalMux t1442 (
    .I(seg_1_22_sp4_h_r_9_9971),
    .O(seg_1_22_local_g1_1_9851)
  );
  Span4Mux_h0 t1443 (
    .I(seg_1_22_sp4_v_t_44_5095),
    .O(seg_1_22_sp4_h_r_9_9971)
  );
  LocalMux t1444 (
    .I(seg_1_22_sp4_h_r_14_4852),
    .O(seg_1_22_local_g0_6_9848)
  );
  Span4Mux_h1 t1445 (
    .I(seg_0_22_sp4_v_t_47_4900),
    .O(seg_1_22_sp4_h_r_14_4852)
  );
  LocalMux t1446 (
    .I(seg_1_1_lutff_2_out_103),
    .O(seg_1_1_local_g0_2_6717)
  );
  LocalMux t1447 (
    .I(seg_1_2_neigh_op_bot_2_103),
    .O(seg_1_2_local_g1_2_6912)
  );
  LocalMux t1448 (
    .I(seg_1_1_lutff_5_out_106),
    .O(seg_1_1_local_g0_5_6720)
  );
  LocalMux t1449 (
    .I(seg_1_2_neigh_op_bot_5_106),
    .O(seg_1_2_local_g1_5_6915)
  );
  CascadeMux t145 (
    .I(net_15179),
    .O(net_15179_cascademuxed)
  );
  LocalMux t1450 (
    .I(seg_1_1_lutff_6_out_107),
    .O(seg_1_1_local_g3_6_6745)
  );
  LocalMux t1451 (
    .I(seg_1_1_lutff_7_out_108),
    .O(seg_1_1_local_g1_7_6730)
  );
  LocalMux t1452 (
    .I(seg_2_3_sp4_v_b_5_6871),
    .O(seg_2_3_local_g0_5_11562)
  );
  LocalMux t1453 (
    .I(seg_1_3_sp4_r_v_b_21_6889),
    .O(seg_1_3_local_g3_5_7078)
  );
  LocalMux t1454 (
    .I(seg_6_4_sp4_h_r_8_27023),
    .O(seg_6_4_local_g0_0_26939)
  );
  Span4Mux_h0 t1455 (
    .I(seg_6_4_sp4_h_l_45_11784),
    .O(seg_6_4_sp4_h_r_8_27023)
  );
  Span4Mux_h4 t1456 (
    .I(seg_2_4_sp4_v_b_8_6889),
    .O(seg_6_4_sp4_h_l_45_11784)
  );
  LocalMux t1457 (
    .I(seg_1_4_sp4_v_b_11_292),
    .O(seg_1_4_local_g0_3_7199)
  );
  LocalMux t1458 (
    .I(seg_2_2_neigh_op_lft_1_117),
    .O(seg_2_2_local_g0_1_11435)
  );
  LocalMux t1459 (
    .I(seg_2_2_neigh_op_lft_2_118),
    .O(seg_2_2_local_g0_2_11436)
  );
  LocalMux t1460 (
    .I(seg_1_1_neigh_op_top_3_119),
    .O(seg_1_1_local_g1_3_6726)
  );
  LocalMux t1461 (
    .I(seg_1_2_lutff_3_out_119),
    .O(seg_1_2_local_g0_3_6905)
  );
  LocalMux t1462 (
    .I(seg_1_2_lutff_4_out_120),
    .O(seg_1_2_local_g2_4_6922)
  );
  LocalMux t1463 (
    .I(seg_2_2_neigh_op_lft_4_120),
    .O(seg_2_2_local_g0_4_11438)
  );
  LocalMux t1464 (
    .I(seg_1_3_neigh_op_bot_5_121),
    .O(seg_1_3_local_g1_5_7062)
  );
  LocalMux t1465 (
    .I(seg_2_2_neigh_op_lft_5_121),
    .O(seg_2_2_local_g1_5_11447)
  );
  LocalMux t1466 (
    .I(seg_1_1_neigh_op_top_6_122),
    .O(seg_1_1_local_g0_6_6721)
  );
  LocalMux t1467 (
    .I(seg_2_1_neigh_op_tnl_7_123),
    .O(seg_2_1_local_g3_7_11302)
  );
  LocalMux t1468 (
    .I(seg_2_2_sp4_h_r_41_523),
    .O(seg_2_2_local_g2_1_11451)
  );
  LocalMux t1469 (
    .I(seg_1_3_lutff_0_out_451),
    .O(seg_1_3_local_g2_0_7065)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t147 (
    .carryinitin(),
    .carryinitout(t146)
  );
  LocalMux t1470 (
    .I(seg_1_4_neigh_op_bot_0_451),
    .O(seg_1_4_local_g0_0_7196)
  );
  LocalMux t1471 (
    .I(seg_1_3_lutff_1_out_452),
    .O(seg_1_3_local_g1_1_7058)
  );
  LocalMux t1472 (
    .I(seg_1_4_neigh_op_bot_1_452),
    .O(seg_1_4_local_g1_1_7205)
  );
  LocalMux t1473 (
    .I(seg_1_2_neigh_op_top_2_453),
    .O(seg_1_2_local_g0_2_6904)
  );
  LocalMux t1474 (
    .I(seg_1_3_lutff_2_out_453),
    .O(seg_1_3_local_g3_2_7075)
  );
  LocalMux t1475 (
    .I(seg_2_3_neigh_op_lft_2_453),
    .O(seg_2_3_local_g1_2_11567)
  );
  LocalMux t1476 (
    .I(seg_1_3_lutff_3_out_454),
    .O(seg_1_3_local_g0_3_7052)
  );
  LocalMux t1477 (
    .I(seg_1_4_neigh_op_bot_3_454),
    .O(seg_1_4_local_g1_3_7207)
  );
  LocalMux t1478 (
    .I(seg_2_4_neigh_op_bnl_3_454),
    .O(seg_2_4_local_g2_3_11699)
  );
  LocalMux t1479 (
    .I(seg_1_3_lutff_4_out_455),
    .O(seg_1_3_local_g3_4_7077)
  );
  CascadeMux t148 (
    .I(net_15300),
    .O(net_15300_cascademuxed)
  );
  LocalMux t1480 (
    .I(seg_2_2_neigh_op_tnl_4_455),
    .O(seg_2_2_local_g2_4_11454)
  );
  LocalMux t1481 (
    .I(seg_2_3_neigh_op_lft_4_455),
    .O(seg_2_3_local_g0_4_11561)
  );
  LocalMux t1482 (
    .I(seg_1_2_neigh_op_top_5_456),
    .O(seg_1_2_local_g0_5_6907)
  );
  LocalMux t1483 (
    .I(seg_2_4_neigh_op_bnl_5_456),
    .O(seg_2_4_local_g3_5_11709)
  );
  LocalMux t1484 (
    .I(seg_2_4_neigh_op_bnl_6_457),
    .O(seg_2_4_local_g3_6_11710)
  );
  LocalMux t1485 (
    .I(seg_1_2_neigh_op_top_7_458),
    .O(seg_1_2_local_g0_7_6909)
  );
  LocalMux t1486 (
    .I(seg_1_3_lutff_7_out_458),
    .O(seg_1_3_local_g2_7_7072)
  );
  LocalMux t1487 (
    .I(seg_2_3_sp4_h_r_23_7169),
    .O(seg_2_3_local_g1_7_11572)
  );
  LocalMux t1488 (
    .I(seg_6_3_sp4_h_r_12_23145),
    .O(seg_6_3_local_g1_4_26849)
  );
  Span4Mux_h1 t1489 (
    .I(seg_5_3_sp4_h_l_47_7169),
    .O(seg_6_3_sp4_h_r_12_23145)
  );
  CascadeMux t149 (
    .I(net_15306),
    .O(net_15306_cascademuxed)
  );
  LocalMux t1490 (
    .I(seg_6_3_sp4_h_r_24_19313),
    .O(seg_6_3_local_g2_0_26853)
  );
  Span4Mux_h2 t1491 (
    .I(seg_4_3_sp4_h_l_44_788),
    .O(seg_6_3_sp4_h_r_24_19313)
  );
  LocalMux t1492 (
    .I(seg_6_4_sp4_v_b_38_23281),
    .O(seg_6_4_local_g2_6_26961)
  );
  Span4Mux_v1 t1493 (
    .I(seg_6_3_sp4_h_l_38_11656),
    .O(seg_6_4_sp4_v_b_38_23281)
  );
  Span4Mux_h4 t1494 (
    .I(seg_2_3_sp4_h_l_38_761),
    .O(seg_6_3_sp4_h_l_38_11656)
  );
  LocalMux t1495 (
    .I(seg_6_3_sp4_h_r_21_23154),
    .O(seg_6_3_local_g1_5_26850)
  );
  Span4Mux_h1 t1496 (
    .I(seg_5_3_sp4_h_l_45_7177),
    .O(seg_6_3_sp4_h_r_21_23154)
  );
  LocalMux t1497 (
    .I(seg_1_3_neigh_op_top_1_679),
    .O(seg_1_3_local_g0_1_7050)
  );
  LocalMux t1498 (
    .I(seg_2_4_neigh_op_lft_2_680),
    .O(seg_2_4_local_g1_2_11690)
  );
  LocalMux t1499 (
    .I(seg_2_5_neigh_op_bnl_2_680),
    .O(seg_2_5_local_g2_2_11821)
  );
  CascadeMux t15 (
    .I(net_7096),
    .O(net_7096_cascademuxed)
  );
  CascadeMux t150 (
    .I(net_15312),
    .O(net_15312_cascademuxed)
  );
  LocalMux t1500 (
    .I(seg_1_3_neigh_op_top_3_681),
    .O(seg_1_3_local_g1_3_7060)
  );
  LocalMux t1501 (
    .I(seg_2_4_neigh_op_lft_4_682),
    .O(seg_2_4_local_g0_4_11684)
  );
  LocalMux t1502 (
    .I(seg_1_4_lutff_5_out_683),
    .O(seg_1_4_local_g0_5_7201)
  );
  LocalMux t1503 (
    .I(seg_2_4_neigh_op_lft_5_683),
    .O(seg_2_4_local_g1_5_11693)
  );
  LocalMux t1504 (
    .I(seg_1_4_lutff_6_out_684),
    .O(seg_1_4_local_g2_6_7218)
  );
  LocalMux t1505 (
    .I(seg_1_5_neigh_op_bot_6_684),
    .O(seg_1_5_local_g1_6_7357)
  );
  LocalMux t1506 (
    .I(seg_2_4_neigh_op_lft_7_685),
    .O(seg_2_4_local_g1_7_11695)
  );
  LocalMux t1507 (
    .I(seg_1_5_lutff_0_out_905),
    .O(seg_1_5_local_g2_0_7359)
  );
  LocalMux t1508 (
    .I(seg_1_4_neigh_op_top_5_910),
    .O(seg_1_4_local_g1_5_7209)
  );
  LocalMux t1509 (
    .I(seg_1_5_lutff_5_out_910),
    .O(seg_1_5_local_g2_5_7364)
  );
  CascadeMux t151 (
    .I(net_15318),
    .O(net_15318_cascademuxed)
  );
  LocalMux t1510 (
    .I(seg_2_5_neigh_op_lft_6_911),
    .O(seg_2_5_local_g0_6_11809)
  );
  LocalMux t1511 (
    .I(seg_0_17_sp4_v_b_6_2928),
    .O(seg_0_17_local_g1_6_3594)
  );
  Span4Mux_v4 t1512 (
    .I(seg_0_13_sp4_v_b_3_2090),
    .O(seg_0_17_sp4_v_b_6_2928)
  );
  Span4Mux_v4 t1513 (
    .I(seg_0_9_sp4_v_b_3_1240),
    .O(seg_0_13_sp4_v_b_3_2090)
  );
  Span4Mux_v4 t1514 (
    .I(seg_0_5_sp4_h_r_3_1201),
    .O(seg_0_9_sp4_v_b_3_1240)
  );
  LocalMux t1515 (
    .I(seg_0_17_sp4_v_b_3_2923),
    .O(seg_0_17_local_g0_3_3583)
  );
  Span4Mux_v4 t1516 (
    .I(seg_0_13_sp4_v_b_7_2094),
    .O(seg_0_17_sp4_v_b_3_2923)
  );
  Span4Mux_v4 t1517 (
    .I(seg_0_9_sp4_v_b_7_1244),
    .O(seg_0_13_sp4_v_b_7_2094)
  );
  Span4Mux_v4 t1518 (
    .I(seg_0_5_sp4_h_r_7_1223),
    .O(seg_0_9_sp4_v_b_7_1244)
  );
  LocalMux t1519 (
    .I(seg_4_4_sp4_v_b_14_15373),
    .O(seg_4_4_local_g0_6_19348)
  );
  CascadeMux t152 (
    .I(net_15330),
    .O(net_15330_cascademuxed)
  );
  Span4Mux_v1 t1520 (
    .I(seg_4_5_sp4_h_l_44_1225),
    .O(seg_4_4_sp4_v_b_14_15373)
  );
  LocalMux t1521 (
    .I(seg_0_7_sp4_v_b_35_1248),
    .O(seg_0_7_local_g2_3_1479)
  );
  Span4Mux_v2 t1522 (
    .I(seg_0_5_sp4_h_r_11_1181),
    .O(seg_0_7_sp4_v_b_35_1248)
  );
  LocalMux t1523 (
    .I(seg_0_17_sp4_v_b_5_2925),
    .O(seg_0_17_local_g0_5_3585)
  );
  Span4Mux_v4 t1524 (
    .I(seg_0_13_sp4_v_b_2_2091),
    .O(seg_0_17_sp4_v_b_5_2925)
  );
  Span4Mux_v4 t1525 (
    .I(seg_0_9_sp4_v_b_11_1248),
    .O(seg_0_13_sp4_v_b_2_2091)
  );
  Span4Mux_v4 t1526 (
    .I(seg_0_5_sp4_h_r_11_1181),
    .O(seg_0_9_sp4_v_b_11_1248)
  );
  LocalMux t1527 (
    .I(seg_2_2_sp4_v_b_36_7032),
    .O(seg_2_2_local_g3_4_11462)
  );
  LocalMux t1528 (
    .I(seg_0_7_sp4_h_r_40_1627),
    .O(seg_0_7_local_g2_0_1476)
  );
  Span4Mux_h1 t1529 (
    .I(seg_1_7_sp4_v_b_0_1017),
    .O(seg_0_7_sp4_h_r_40_1627)
  );
  CascadeMux t153 (
    .I(net_15342),
    .O(net_15342_cascademuxed)
  );
  LocalMux t1530 (
    .I(seg_0_7_sp4_h_r_47_1634),
    .O(seg_0_7_local_g2_7_1483)
  );
  Span4Mux_h1 t1531 (
    .I(seg_1_7_sp4_v_b_10_1027),
    .O(seg_0_7_sp4_h_r_47_1634)
  );
  LocalMux t1532 (
    .I(seg_0_7_sp4_r_v_b_22_1236),
    .O(seg_0_7_local_g3_6_1490)
  );
  LocalMux t1533 (
    .I(seg_0_17_sp4_r_v_b_10_3147),
    .O(seg_0_17_local_g2_2_3598)
  );
  Span4Mux_v4 t1534 (
    .I(seg_1_13_sp4_v_b_7_2292),
    .O(seg_0_17_sp4_r_v_b_10_3147)
  );
  Span4Mux_v4 t1535 (
    .I(seg_1_9_sp4_v_b_11_1442),
    .O(seg_1_13_sp4_v_b_7_2292)
  );
  Span4Mux_v4 t1536 (
    .I(seg_1_5_sp4_v_b_8_571),
    .O(seg_1_9_sp4_v_b_11_1442)
  );
  LocalMux t1537 (
    .I(seg_1_6_lutff_1_out_1131),
    .O(seg_1_6_local_g0_1_7491)
  );
  LocalMux t1538 (
    .I(seg_0_7_neigh_op_bnr_3_1133),
    .O(seg_0_7_local_g1_3_1471)
  );
  LocalMux t1539 (
    .I(seg_1_6_lutff_5_out_1135),
    .O(seg_1_6_local_g3_5_7519)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t154 (
    .carryinitin(net_19170),
    .carryinitout(net_19214)
  );
  LocalMux t1540 (
    .I(seg_0_7_neigh_op_bnr_6_1136),
    .O(seg_0_7_local_g1_6_1474)
  );
  LocalMux t1541 (
    .I(seg_0_17_sp4_r_v_b_12_3346),
    .O(seg_0_17_local_g2_4_3600)
  );
  Sp12to4 t1542 (
    .I(seg_1_17_sp12_v_b_1_7459),
    .O(seg_0_17_sp4_r_v_b_12_3346)
  );
  LocalMux t1543 (
    .I(seg_1_8_sp4_v_b_16_1436),
    .O(seg_1_8_local_g1_0_7792)
  );
  LocalMux t1544 (
    .I(seg_0_17_sp4_r_v_b_9_3144),
    .O(seg_0_17_local_g2_1_3597)
  );
  Span4Mux_v4 t1545 (
    .I(seg_1_13_sp4_v_b_9_2294),
    .O(seg_0_17_sp4_r_v_b_9_3144)
  );
  Span4Mux_v4 t1546 (
    .I(seg_1_9_sp4_v_b_9_1440),
    .O(seg_1_13_sp4_v_b_9_2294)
  );
  LocalMux t1547 (
    .I(seg_2_7_neigh_op_lft_1_1337),
    .O(seg_2_7_local_g0_1_12050)
  );
  LocalMux t1548 (
    .I(seg_1_8_lutff_0_out_1544),
    .O(seg_1_8_local_g3_0_7808)
  );
  LocalMux t1549 (
    .I(seg_1_8_lutff_1_out_1545),
    .O(seg_1_8_local_g2_1_7801)
  );
  CascadeMux t155 (
    .I(net_15423),
    .O(net_15423_cascademuxed)
  );
  LocalMux t1550 (
    .I(seg_1_8_lutff_2_out_1546),
    .O(seg_1_8_local_g2_2_7802)
  );
  LocalMux t1551 (
    .I(seg_0_7_neigh_op_tnr_3_1547),
    .O(seg_0_7_local_g3_3_1487)
  );
  LocalMux t1552 (
    .I(seg_0_7_neigh_op_tnr_4_1548),
    .O(seg_0_7_local_g3_4_1488)
  );
  LocalMux t1553 (
    .I(seg_1_8_lutff_6_out_1550),
    .O(seg_1_8_local_g1_6_7798)
  );
  LocalMux t1554 (
    .I(seg_0_7_neigh_op_tnr_7_1551),
    .O(seg_0_7_local_g3_7_1491)
  );
  LocalMux t1555 (
    .I(seg_9_7_sp4_v_b_23_34275),
    .O(seg_9_7_local_g0_7_38242)
  );
  Span4Mux_v1 t1556 (
    .I(seg_9_8_sp4_h_l_47_23761),
    .O(seg_9_7_sp4_v_b_23_34275)
  );
  Span4Mux_h4 t1557 (
    .I(seg_5_8_sp4_h_l_47_7904),
    .O(seg_9_8_sp4_h_l_47_23761)
  );
  LocalMux t1558 (
    .I(seg_0_17_sp4_r_v_b_23_3357),
    .O(seg_0_17_local_g3_7_3611)
  );
  Span4Mux_v3 t1559 (
    .I(seg_1_14_sp4_v_b_2_2495),
    .O(seg_0_17_sp4_r_v_b_23_3357)
  );
  CascadeMux t156 (
    .I(net_15429),
    .O(net_15429_cascademuxed)
  );
  Span4Mux_v4 t1560 (
    .I(seg_1_10_sp4_v_b_6_1647),
    .O(seg_1_14_sp4_v_b_2_2495)
  );
  LocalMux t1561 (
    .I(seg_0_17_sp4_r_v_b_31_3558),
    .O(seg_0_17_local_g1_7_3595)
  );
  Span4Mux_v2 t1562 (
    .I(seg_1_15_sp4_v_b_11_2710),
    .O(seg_0_17_sp4_r_v_b_31_3558)
  );
  Span4Mux_v4 t1563 (
    .I(seg_1_11_sp4_v_b_3_1851),
    .O(seg_1_15_sp4_v_b_11_2710)
  );
  LocalMux t1564 (
    .I(seg_0_17_sp4_r_v_b_28_3557),
    .O(seg_0_17_local_g1_4_3592)
  );
  Span4Mux_v2 t1565 (
    .I(seg_1_15_sp4_v_b_8_2709),
    .O(seg_0_17_sp4_r_v_b_28_3557)
  );
  Span4Mux_v4 t1566 (
    .I(seg_1_11_sp4_v_b_5_1853),
    .O(seg_1_15_sp4_v_b_8_2709)
  );
  LocalMux t1567 (
    .I(seg_2_9_neigh_op_lft_5_1758),
    .O(seg_2_9_local_g0_5_12300)
  );
  LocalMux t1568 (
    .I(seg_2_9_neigh_op_lft_7_1760),
    .O(seg_2_9_local_g0_7_12302)
  );
  LocalMux t1569 (
    .I(seg_0_16_sp4_v_b_22_2931),
    .O(seg_0_16_local_g0_6_3380)
  );
  CascadeMux t157 (
    .I(net_15441),
    .O(net_15441_cascademuxed)
  );
  Span4Mux_v3 t1570 (
    .I(seg_0_13_sp4_v_b_11_2098),
    .O(seg_0_16_sp4_v_b_22_2931)
  );
  Span4Mux_v4 t1571 (
    .I(seg_0_9_sp4_h_r_5_2071),
    .O(seg_0_13_sp4_v_b_11_2098)
  );
  LocalMux t1572 (
    .I(seg_0_11_sp4_h_r_34_2472),
    .O(seg_0_11_local_g2_2_2332)
  );
  Span4Mux_h2 t1573 (
    .I(seg_2_11_sp4_v_b_5_7918),
    .O(seg_0_11_sp4_h_r_34_2472)
  );
  LocalMux t1574 (
    .I(seg_0_16_sp4_h_r_31_3529),
    .O(seg_0_16_local_g2_7_3397)
  );
  Span4Mux_h2 t1575 (
    .I(seg_2_16_sp4_v_b_7_8655),
    .O(seg_0_16_sp4_h_r_31_3529)
  );
  Span4Mux_v4 t1576 (
    .I(seg_2_12_sp4_v_b_4_8066),
    .O(seg_2_16_sp4_v_b_7_8655)
  );
  LocalMux t1577 (
    .I(seg_0_16_sp4_h_r_33_3531),
    .O(seg_0_16_local_g3_1_3399)
  );
  Span4Mux_h2 t1578 (
    .I(seg_2_16_sp4_v_b_4_8654),
    .O(seg_0_16_sp4_h_r_33_3531)
  );
  Span4Mux_v4 t1579 (
    .I(seg_2_12_sp4_v_b_8_8070),
    .O(seg_2_16_sp4_v_b_4_8654)
  );
  CascadeMux t158 (
    .I(net_15447),
    .O(net_15447_cascademuxed)
  );
  LocalMux t1580 (
    .I(seg_0_11_sp4_r_v_b_0_1850),
    .O(seg_0_11_local_g1_0_2322)
  );
  LocalMux t1581 (
    .I(seg_0_11_sp4_r_v_b_8_1858),
    .O(seg_0_11_local_g2_0_2330)
  );
  LocalMux t1582 (
    .I(seg_0_11_sp4_h_r_47_2486),
    .O(seg_0_11_local_g2_7_2337)
  );
  Span4Mux_h1 t1583 (
    .I(seg_1_11_sp4_v_b_10_1860),
    .O(seg_0_11_sp4_h_r_47_2486)
  );
  LocalMux t1584 (
    .I(seg_0_16_sp4_r_v_b_44_3560),
    .O(seg_0_16_local_g3_4_3402)
  );
  Span4Mux_v1 t1585 (
    .I(seg_1_15_sp4_v_b_6_2707),
    .O(seg_0_16_sp4_r_v_b_44_3560)
  );
  Span4Mux_v4 t1586 (
    .I(seg_1_11_sp4_v_b_10_1860),
    .O(seg_1_15_sp4_v_b_6_2707)
  );
  LocalMux t1587 (
    .I(seg_0_11_sp4_r_v_b_12_2076),
    .O(seg_0_11_local_g2_4_2334)
  );
  LocalMux t1588 (
    .I(seg_0_16_sp4_r_v_b_1_2909),
    .O(seg_0_16_local_g1_1_3383)
  );
  Span4Mux_v4 t1589 (
    .I(seg_1_12_sp4_v_b_1_2076),
    .O(seg_0_16_sp4_r_v_b_1_2909)
  );
  CascadeMux t159 (
    .I(net_15453),
    .O(net_15453_cascademuxed)
  );
  LocalMux t1590 (
    .I(seg_0_11_sp4_r_v_b_20_2084),
    .O(seg_0_11_local_g3_4_2342)
  );
  Span4Mux_v1 t1591 (
    .I(seg_1_12_sp4_h_l_38_2684),
    .O(seg_0_11_sp4_r_v_b_20_2084)
  );
  Span4Mux_h0 t1592 (
    .I(seg_1_12_sp4_v_b_3_2078),
    .O(seg_1_12_sp4_h_l_38_2684)
  );
  LocalMux t1593 (
    .I(seg_0_16_sp4_r_v_b_6_2916),
    .O(seg_0_16_local_g1_6_3388)
  );
  Span4Mux_v4 t1594 (
    .I(seg_1_12_sp4_v_b_3_2078),
    .O(seg_0_16_sp4_r_v_b_6_2916)
  );
  LocalMux t1595 (
    .I(seg_1_9_neigh_op_top_0_1965),
    .O(seg_1_9_local_g0_0_7931)
  );
  LocalMux t1596 (
    .I(seg_2_9_neigh_op_tnl_1_1966),
    .O(seg_2_9_local_g2_1_12312)
  );
  LocalMux t1597 (
    .I(seg_1_10_lutff_3_out_1968),
    .O(seg_1_10_local_g0_3_8081)
  );
  LocalMux t1598 (
    .I(seg_1_10_lutff_4_out_1969),
    .O(seg_1_10_local_g2_4_8098)
  );
  LocalMux t1599 (
    .I(seg_1_10_lutff_5_out_1970),
    .O(seg_1_10_local_g0_5_8083)
  );
  CascadeMux t16 (
    .I(net_7108),
    .O(net_7108_cascademuxed)
  );
  CascadeMux t160 (
    .I(net_15459),
    .O(net_15459_cascademuxed)
  );
  LocalMux t1600 (
    .I(seg_2_10_neigh_op_lft_6_1971),
    .O(seg_2_10_local_g1_6_12432)
  );
  LocalMux t1601 (
    .I(seg_1_10_lutff_7_out_1972),
    .O(seg_1_10_local_g0_7_8085)
  );
  LocalMux t1602 (
    .I(seg_16_10_sp4_h_r_10_65515),
    .O(seg_16_10_local_g0_2_65421)
  );
  Span4Mux_h0 t1603 (
    .I(seg_16_10_sp4_h_l_47_50193),
    .O(seg_16_10_sp4_h_r_10_65515)
  );
  Span4Mux_h4 t1604 (
    .I(seg_12_10_sp4_h_l_42_34876),
    .O(seg_16_10_sp4_h_l_47_50193)
  );
  Span4Mux_h4 t1605 (
    .I(seg_8_10_sp4_h_l_41_20180),
    .O(seg_12_10_sp4_h_l_42_34876)
  );
  Span4Mux_h4 t1606 (
    .I(seg_4_10_sp4_h_l_36_2239),
    .O(seg_8_10_sp4_h_l_41_20180)
  );
  LocalMux t1607 (
    .I(seg_5_7_sp4_v_b_41_19822),
    .O(seg_5_7_local_g3_1_23567)
  );
  Span4Mux_v3 t1608 (
    .I(seg_5_10_sp4_h_l_41_8202),
    .O(seg_5_7_sp4_v_b_41_19822)
  );
  LocalMux t1609 (
    .I(seg_5_10_sp4_h_r_7_24014),
    .O(seg_5_10_local_g0_7_23918)
  );
  CascadeMux t161 (
    .I(net_15465),
    .O(net_15465_cascademuxed)
  );
  Span4Mux_h0 t1610 (
    .I(seg_5_10_sp4_h_l_41_8202),
    .O(seg_5_10_sp4_h_r_7_24014)
  );
  LocalMux t1611 (
    .I(seg_16_10_sp4_h_r_36_54023),
    .O(seg_16_10_local_g2_4_65439)
  );
  Span4Mux_h3 t1612 (
    .I(seg_13_10_sp4_h_l_47_38700),
    .O(seg_16_10_sp4_h_r_36_54023)
  );
  Span4Mux_h4 t1613 (
    .I(seg_9_10_sp4_h_l_42_24014),
    .O(seg_13_10_sp4_h_l_47_38700)
  );
  Span4Mux_h4 t1614 (
    .I(seg_5_10_sp4_h_l_41_8202),
    .O(seg_9_10_sp4_h_l_42_24014)
  );
  LocalMux t1615 (
    .I(seg_2_7_sp4_h_r_5_12150),
    .O(seg_2_7_local_g0_5_12054)
  );
  Span4Mux_h0 t1616 (
    .I(seg_2_7_sp4_v_t_37_7915),
    .O(seg_2_7_sp4_h_r_5_12150)
  );
  LocalMux t1617 (
    .I(seg_2_8_sp4_v_b_37_7915),
    .O(seg_2_8_local_g2_5_12193)
  );
  LocalMux t1618 (
    .I(seg_3_8_sp4_h_r_16_12273),
    .O(seg_3_8_local_g0_0_16003)
  );
  Span4Mux_h1 t1619 (
    .I(seg_2_8_sp4_v_t_40_8065),
    .O(seg_3_8_sp4_h_r_16_12273)
  );
  CascadeMux t162 (
    .I(net_15546),
    .O(net_15546_cascademuxed)
  );
  LocalMux t1620 (
    .I(seg_2_7_sp4_v_b_40_7771),
    .O(seg_2_7_local_g2_0_12065)
  );
  LocalMux t1621 (
    .I(seg_2_8_sp4_v_b_29_7771),
    .O(seg_2_8_local_g3_5_12201)
  );
  LocalMux t1622 (
    .I(seg_2_10_neigh_op_tnl_0_2190),
    .O(seg_2_10_local_g3_0_12442)
  );
  LocalMux t1623 (
    .I(seg_2_10_neigh_op_tnl_1_2191),
    .O(seg_2_10_local_g3_1_12443)
  );
  LocalMux t1624 (
    .I(seg_1_11_lutff_2_out_2192),
    .O(seg_1_11_local_g1_2_8235)
  );
  LocalMux t1625 (
    .I(seg_2_10_neigh_op_tnl_4_2194),
    .O(seg_2_10_local_g3_4_12446)
  );
  LocalMux t1626 (
    .I(seg_2_10_neigh_op_tnl_5_2195),
    .O(seg_2_10_local_g2_5_12439)
  );
  LocalMux t1627 (
    .I(seg_1_11_lutff_7_out_2197),
    .O(seg_1_11_local_g0_7_8232)
  );
  LocalMux t1628 (
    .I(seg_5_10_sp4_v_b_19_19947),
    .O(seg_5_10_local_g0_3_23914)
  );
  Span4Mux_v1 t1629 (
    .I(seg_5_11_sp4_h_l_43_8351),
    .O(seg_5_10_sp4_v_b_19_19947)
  );
  CascadeMux t163 (
    .I(net_15564),
    .O(net_15564_cascademuxed)
  );
  LocalMux t1630 (
    .I(seg_12_10_sp4_r_v_b_17_49962),
    .O(seg_12_10_local_g3_1_50122)
  );
  Span4Mux_v1 t1631 (
    .I(seg_13_11_sp4_h_l_47_38823),
    .O(seg_12_10_sp4_r_v_b_17_49962)
  );
  Span4Mux_h4 t1632 (
    .I(seg_9_11_sp4_h_l_39_24132),
    .O(seg_13_11_sp4_h_l_47_38823)
  );
  Span4Mux_h4 t1633 (
    .I(seg_5_11_sp4_h_l_43_8351),
    .O(seg_9_11_sp4_h_l_39_24132)
  );
  LocalMux t1634 (
    .I(seg_4_12_sp4_h_r_34_12760),
    .O(seg_4_12_local_g3_2_20352)
  );
  Span4Mux_h2 t1635 (
    .I(seg_2_12_sp4_v_b_10_8072),
    .O(seg_4_12_sp4_h_r_34_12760)
  );
  LocalMux t1636 (
    .I(seg_2_7_sp4_h_r_7_12152),
    .O(seg_2_7_local_g0_7_12056)
  );
  Span4Mux_h0 t1637 (
    .I(seg_2_7_sp4_v_t_42_7920),
    .O(seg_2_7_sp4_h_r_7_12152)
  );
  LocalMux t1638 (
    .I(seg_0_6_sp4_r_v_b_42_1438),
    .O(seg_0_6_local_g3_2_1280)
  );
  Span4Mux_v3 t1639 (
    .I(seg_1_9_sp4_v_t_41_2291),
    .O(seg_0_6_sp4_r_v_b_42_1438)
  );
  CascadeMux t164 (
    .I(net_15570),
    .O(net_15570_cascademuxed)
  );
  LocalMux t1640 (
    .I(seg_0_24_sp4_r_v_b_18_4883),
    .O(seg_0_24_local_g3_2_5141)
  );
  Span4Mux_v3 t1641 (
    .I(seg_1_21_sp4_v_b_4_3974),
    .O(seg_0_24_sp4_r_v_b_18_4883)
  );
  Span4Mux_v4 t1642 (
    .I(seg_1_17_sp4_v_b_4_3141),
    .O(seg_1_21_sp4_v_b_4_3974)
  );
  Span4Mux_v4 t1643 (
    .I(seg_1_13_sp4_v_b_4_2291),
    .O(seg_1_17_sp4_v_b_4_3141)
  );
  LocalMux t1644 (
    .I(seg_1_7_sp4_h_r_6_7763),
    .O(seg_1_7_local_g1_6_7651)
  );
  Span4Mux_h0 t1645 (
    .I(seg_1_7_sp4_v_t_43_1856),
    .O(seg_1_7_sp4_h_r_6_7763)
  );
  LocalMux t1646 (
    .I(seg_1_12_lutff_3_out_2399),
    .O(seg_1_12_local_g0_3_8375)
  );
  LocalMux t1647 (
    .I(seg_1_12_lutff_5_out_2401),
    .O(seg_1_12_local_g0_5_8377)
  );
  LocalMux t1648 (
    .I(seg_1_12_lutff_6_out_2402),
    .O(seg_1_12_local_g0_6_8378)
  );
  LocalMux t1649 (
    .I(seg_3_12_sp4_h_r_3_16594),
    .O(seg_3_12_local_g0_3_16498)
  );
  CascadeMux t165 (
    .I(net_15705),
    .O(net_15705_cascademuxed)
  );
  Span4Mux_h0 t1650 (
    .I(seg_3_12_sp4_h_l_37_2657),
    .O(seg_3_12_sp4_h_r_3_16594)
  );
  LocalMux t1651 (
    .I(seg_3_12_sp4_h_r_12_12759),
    .O(seg_3_12_local_g1_4_16507)
  );
  Span4Mux_h1 t1652 (
    .I(seg_2_12_sp4_h_l_36_2670),
    .O(seg_3_12_sp4_h_r_12_12759)
  );
  LocalMux t1653 (
    .I(seg_3_10_sp4_h_r_13_12512),
    .O(seg_3_10_local_g0_5_16254)
  );
  Span4Mux_h1 t1654 (
    .I(seg_2_10_sp4_v_t_42_8361),
    .O(seg_3_10_sp4_h_r_13_12512)
  );
  LocalMux t1655 (
    .I(seg_3_10_sp4_h_r_20_12523),
    .O(seg_3_10_local_g1_4_16261)
  );
  Span4Mux_h1 t1656 (
    .I(seg_2_10_sp4_v_t_44_8363),
    .O(seg_3_10_sp4_h_r_20_12523)
  );
  LocalMux t1657 (
    .I(seg_4_13_sp4_h_r_37_8637),
    .O(seg_4_13_local_g2_5_20470)
  );
  LocalMux t1658 (
    .I(seg_4_13_sp4_h_r_39_8641),
    .O(seg_4_13_local_g2_7_20472)
  );
  LocalMux t1659 (
    .I(seg_4_13_sp4_h_r_11_20546),
    .O(seg_4_13_local_g0_3_20452)
  );
  CascadeMux t166 (
    .I(net_15816),
    .O(net_15816_cascademuxed)
  );
  Span4Mux_h0 t1660 (
    .I(seg_4_13_sp4_h_l_46_2864),
    .O(seg_4_13_sp4_h_r_11_20546)
  );
  LocalMux t1661 (
    .I(seg_4_13_sp4_h_r_16_16719),
    .O(seg_4_13_local_g0_0_20449)
  );
  Span4Mux_h1 t1662 (
    .I(seg_3_13_sp4_h_l_39_2868),
    .O(seg_4_13_sp4_h_r_16_16719)
  );
  LocalMux t1663 (
    .I(seg_4_13_sp4_h_r_17_16718),
    .O(seg_4_13_local_g0_1_20450)
  );
  Span4Mux_h1 t1664 (
    .I(seg_3_13_sp4_h_l_41_2870),
    .O(seg_4_13_sp4_h_r_17_16718)
  );
  LocalMux t1665 (
    .I(seg_4_13_sp4_h_r_19_16720),
    .O(seg_4_13_local_g1_3_20460)
  );
  Span4Mux_h1 t1666 (
    .I(seg_3_13_sp4_h_l_43_2872),
    .O(seg_4_13_sp4_h_r_19_16720)
  );
  LocalMux t1667 (
    .I(seg_4_13_sp4_h_r_41_8643),
    .O(seg_4_13_local_g2_1_20466)
  );
  LocalMux t1668 (
    .I(seg_4_13_sp4_h_r_45_8647),
    .O(seg_4_13_local_g3_5_20478)
  );
  LocalMux t1669 (
    .I(seg_2_13_neigh_op_tnl_1_2814),
    .O(seg_2_13_local_g2_1_12804)
  );
  CascadeMux t167 (
    .I(net_15828),
    .O(net_15828_cascademuxed)
  );
  LocalMux t1670 (
    .I(seg_2_13_neigh_op_tnl_3_2816),
    .O(seg_2_13_local_g3_3_12814)
  );
  LocalMux t1671 (
    .I(seg_1_14_lutff_4_out_2817),
    .O(seg_1_14_local_g0_4_8670)
  );
  LocalMux t1672 (
    .I(seg_2_15_neigh_op_bnl_6_2819),
    .O(seg_2_15_local_g3_6_13063)
  );
  LocalMux t1673 (
    .I(seg_1_11_sp4_h_r_45_2470),
    .O(seg_1_11_local_g3_5_8254)
  );
  Span4Mux_h1 t1674 (
    .I(seg_2_11_sp4_v_t_39_8505),
    .O(seg_1_11_sp4_h_r_45_2470)
  );
  LocalMux t1675 (
    .I(seg_1_11_sp4_v_b_37_2493),
    .O(seg_1_11_local_g2_5_8246)
  );
  LocalMux t1676 (
    .I(seg_1_11_sp4_v_b_47_2503),
    .O(seg_1_11_local_g2_7_8248)
  );
  LocalMux t1677 (
    .I(seg_1_12_sp4_v_b_28_2497),
    .O(seg_1_12_local_g2_4_8392)
  );
  LocalMux t1678 (
    .I(seg_1_15_lutff_0_out_3025),
    .O(seg_1_15_local_g0_0_8813)
  );
  LocalMux t1679 (
    .I(seg_1_15_lutff_1_out_3026),
    .O(seg_1_15_local_g3_1_8838)
  );
  CascadeMux t168 (
    .I(net_15915),
    .O(net_15915_cascademuxed)
  );
  LocalMux t1680 (
    .I(seg_2_15_neigh_op_lft_2_3027),
    .O(seg_2_15_local_g1_2_13043)
  );
  LocalMux t1681 (
    .I(seg_1_14_neigh_op_top_3_3028),
    .O(seg_1_14_local_g0_3_8669)
  );
  LocalMux t1682 (
    .I(seg_1_15_lutff_4_out_3029),
    .O(seg_1_15_local_g3_4_8841)
  );
  LocalMux t1683 (
    .I(seg_1_14_neigh_op_top_5_3030),
    .O(seg_1_14_local_g0_5_8671)
  );
  LocalMux t1684 (
    .I(seg_1_15_lutff_6_out_3031),
    .O(seg_1_15_local_g1_6_8827)
  );
  LocalMux t1685 (
    .I(seg_1_14_neigh_op_top_7_3032),
    .O(seg_1_14_local_g0_7_8673)
  );
  LocalMux t1686 (
    .I(seg_1_16_lutff_0_out_3250),
    .O(seg_1_16_local_g3_0_8984)
  );
  LocalMux t1687 (
    .I(seg_2_16_neigh_op_lft_2_3252),
    .O(seg_2_16_local_g0_2_13158)
  );
  LocalMux t1688 (
    .I(seg_2_15_neigh_op_tnl_3_3253),
    .O(seg_2_15_local_g3_3_13060)
  );
  LocalMux t1689 (
    .I(seg_1_16_lutff_4_out_3254),
    .O(seg_1_16_local_g3_4_8988)
  );
  CascadeMux t169 (
    .I(net_15921),
    .O(net_15921_cascademuxed)
  );
  LocalMux t1690 (
    .I(seg_1_16_lutff_5_out_3255),
    .O(seg_1_16_local_g0_5_8965)
  );
  LocalMux t1691 (
    .I(seg_1_16_lutff_6_out_3256),
    .O(seg_1_16_local_g2_6_8982)
  );
  LocalMux t1692 (
    .I(seg_4_16_sp4_h_r_39_9082),
    .O(seg_4_16_local_g2_7_20841)
  );
  LocalMux t1693 (
    .I(seg_2_16_neigh_op_tnl_1_3457),
    .O(seg_2_16_local_g2_1_13173)
  );
  LocalMux t1694 (
    .I(seg_2_16_neigh_op_tnl_2_3458),
    .O(seg_2_16_local_g2_2_13174)
  );
  LocalMux t1695 (
    .I(seg_1_11_sp4_r_v_b_27_8210),
    .O(seg_1_11_local_g0_3_8228)
  );
  Span4Mux_v2 t1696 (
    .I(seg_2_13_sp4_v_t_42_8802),
    .O(seg_1_11_sp4_r_v_b_27_8210)
  );
  LocalMux t1697 (
    .I(seg_1_10_sp4_h_r_11_8199),
    .O(seg_1_10_local_g1_3_8089)
  );
  Span4Mux_h0 t1698 (
    .I(seg_1_10_sp4_v_t_43_2499),
    .O(seg_1_10_sp4_h_r_11_8199)
  );
  Span4Mux_v4 t1699 (
    .I(seg_1_14_sp4_v_t_38_3348),
    .O(seg_1_10_sp4_v_t_43_2499)
  );
  CascadeMux t17 (
    .I(net_7114),
    .O(net_7114_cascademuxed)
  );
  CascadeMux t170 (
    .I(net_15927),
    .O(net_15927_cascademuxed)
  );
  LocalMux t1700 (
    .I(seg_1_17_neigh_op_top_0_3664),
    .O(seg_1_17_local_g0_0_9107)
  );
  LocalMux t1701 (
    .I(seg_1_17_neigh_op_top_1_3665),
    .O(seg_1_17_local_g0_1_9108)
  );
  LocalMux t1702 (
    .I(seg_1_17_neigh_op_top_4_3668),
    .O(seg_1_17_local_g0_4_9111)
  );
  LocalMux t1703 (
    .I(seg_2_17_neigh_op_tnl_6_3670),
    .O(seg_2_17_local_g2_6_13301)
  );
  LocalMux t1704 (
    .I(seg_2_19_neigh_op_lft_0_3873),
    .O(seg_2_19_local_g1_0_13533)
  );
  LocalMux t1705 (
    .I(seg_1_18_neigh_op_top_5_3878),
    .O(seg_1_18_local_g1_5_9267)
  );
  LocalMux t1706 (
    .I(seg_1_18_neigh_op_top_7_3880),
    .O(seg_1_18_local_g0_7_9261)
  );
  LocalMux t1707 (
    .I(seg_1_19_neigh_op_top_1_4086),
    .O(seg_1_19_local_g0_1_9402)
  );
  LocalMux t1708 (
    .I(seg_2_20_neigh_op_lft_2_4087),
    .O(seg_2_20_local_g0_2_13650)
  );
  LocalMux t1709 (
    .I(seg_1_19_neigh_op_top_6_4091),
    .O(seg_1_19_local_g0_6_9407)
  );
  CascadeMux t171 (
    .I(net_15933),
    .O(net_15933_cascademuxed)
  );
  LocalMux t1710 (
    .I(seg_1_19_neigh_op_top_7_4092),
    .O(seg_1_19_local_g1_7_9416)
  );
  LocalMux t1711 (
    .I(seg_2_20_neigh_op_tnl_0_4312),
    .O(seg_2_20_local_g3_0_13672)
  );
  LocalMux t1712 (
    .I(seg_1_18_sp4_v_b_43_3976),
    .O(seg_1_18_local_g3_3_9281)
  );
  LocalMux t1713 (
    .I(seg_1_22_lutff_1_out_4540),
    .O(seg_1_22_local_g0_1_9843)
  );
  LocalMux t1714 (
    .I(seg_1_21_neigh_op_top_5_4544),
    .O(seg_1_21_local_g0_5_9700)
  );
  LocalMux t1715 (
    .I(seg_1_20_sp4_v_b_36_4423),
    .O(seg_1_20_local_g3_4_9576)
  );
  LocalMux t1716 (
    .I(seg_2_22_neigh_op_tnl_2_4768),
    .O(seg_2_22_local_g3_2_13920)
  );
  LocalMux t1717 (
    .I(seg_2_1_lutff_0_out_6673),
    .O(seg_2_1_local_g3_0_11295)
  );
  LocalMux t1718 (
    .I(seg_2_1_lutff_1_out_6674),
    .O(seg_2_1_local_g0_1_11272)
  );
  LocalMux t1719 (
    .I(seg_2_2_neigh_op_bot_3_6676),
    .O(seg_2_2_local_g1_3_11445)
  );
  CascadeMux t172 (
    .I(net_15939),
    .O(net_15939_cascademuxed)
  );
  LocalMux t1720 (
    .I(seg_2_2_neigh_op_bot_5_6678),
    .O(seg_2_2_local_g0_5_11439)
  );
  LocalMux t1721 (
    .I(seg_2_1_lutff_7_out_6680),
    .O(seg_2_1_local_g0_7_11278)
  );
  LocalMux t1722 (
    .I(seg_1_2_sp4_r_v_b_31_6886),
    .O(seg_1_2_local_g1_7_6917)
  );
  LocalMux t1723 (
    .I(seg_1_3_neigh_op_bnr_0_6825),
    .O(seg_1_3_local_g1_0_7057)
  );
  LocalMux t1724 (
    .I(seg_2_2_lutff_0_out_6825),
    .O(seg_2_2_local_g1_0_11442)
  );
  LocalMux t1725 (
    .I(seg_2_3_neigh_op_bot_0_6825),
    .O(seg_2_3_local_g1_0_11565)
  );
  LocalMux t1726 (
    .I(seg_1_2_neigh_op_rgt_1_6826),
    .O(seg_1_2_local_g2_1_6919)
  );
  LocalMux t1727 (
    .I(seg_2_3_neigh_op_bot_1_6826),
    .O(seg_2_3_local_g0_1_11558)
  );
  LocalMux t1728 (
    .I(seg_2_2_lutff_2_out_6827),
    .O(seg_2_2_local_g2_2_11452)
  );
  LocalMux t1729 (
    .I(seg_3_1_neigh_op_tnl_3_6828),
    .O(seg_3_1_local_g3_3_15129)
  );
  CascadeMux t173 (
    .I(net_15945),
    .O(net_15945_cascademuxed)
  );
  LocalMux t1730 (
    .I(seg_2_1_neigh_op_top_4_6829),
    .O(seg_2_1_local_g1_4_11283)
  );
  LocalMux t1731 (
    .I(seg_2_3_neigh_op_bot_4_6829),
    .O(seg_2_3_local_g1_4_11569)
  );
  LocalMux t1732 (
    .I(seg_2_2_lutff_5_out_6830),
    .O(seg_2_2_local_g2_5_11455)
  );
  LocalMux t1733 (
    .I(seg_1_2_neigh_op_rgt_6_6831),
    .O(seg_1_2_local_g2_6_6924)
  );
  LocalMux t1734 (
    .I(seg_2_3_neigh_op_bot_6_6831),
    .O(seg_2_3_local_g0_6_11563)
  );
  LocalMux t1735 (
    .I(seg_1_2_neigh_op_rgt_7_6832),
    .O(seg_1_2_local_g2_7_6925)
  );
  LocalMux t1736 (
    .I(seg_2_2_lutff_7_out_6832),
    .O(seg_2_2_local_g1_7_11449)
  );
  LocalMux t1737 (
    .I(seg_6_4_sp4_v_b_29_23160),
    .O(seg_6_4_local_g3_5_26968)
  );
  Span4Mux_v2 t1738 (
    .I(seg_6_2_sp4_h_l_37_11528),
    .O(seg_6_4_sp4_v_b_29_23160)
  );
  LocalMux t1739 (
    .I(seg_4_1_sp4_r_v_b_22_19058),
    .O(seg_4_1_local_g3_6_18963)
  );
  CascadeMux t174 (
    .I(net_15957),
    .O(net_15957_cascademuxed)
  );
  Span4Mux_v1 t1740 (
    .I(seg_5_2_sp4_h_l_46_7023),
    .O(seg_4_1_sp4_r_v_b_22_19058)
  );
  LocalMux t1741 (
    .I(seg_4_4_sp4_r_v_b_28_19330),
    .O(seg_4_4_local_g0_4_19346)
  );
  Span4Mux_v2 t1742 (
    .I(seg_5_2_sp4_h_l_46_7023),
    .O(seg_4_4_sp4_r_v_b_28_19330)
  );
  LocalMux t1743 (
    .I(seg_5_1_sp4_r_v_b_13_22879),
    .O(seg_5_1_local_g2_5_22785)
  );
  Span4Mux_v1 t1744 (
    .I(seg_6_2_sp4_h_l_43_11536),
    .O(seg_5_1_sp4_r_v_b_13_22879)
  );
  LocalMux t1745 (
    .I(seg_6_4_sp4_v_b_25_23156),
    .O(seg_6_4_local_g2_1_26956)
  );
  Span4Mux_v2 t1746 (
    .I(seg_6_2_sp4_h_l_45_11538),
    .O(seg_6_4_sp4_v_b_25_23156)
  );
  LocalMux t1747 (
    .I(seg_3_4_sp4_v_b_15_11543),
    .O(seg_3_4_local_g1_7_15526)
  );
  LocalMux t1748 (
    .I(seg_2_4_sp4_v_b_16_7036),
    .O(seg_2_4_local_g0_0_11680)
  );
  LocalMux t1749 (
    .I(seg_2_3_lutff_0_out_7008),
    .O(seg_2_3_local_g2_0_11573)
  );
  LocalMux t1750 (
    .I(seg_3_4_neigh_op_bnl_1_7009),
    .O(seg_3_4_local_g3_1_15536)
  );
  LocalMux t1751 (
    .I(seg_2_2_neigh_op_top_2_7010),
    .O(seg_2_2_local_g1_2_11444)
  );
  LocalMux t1752 (
    .I(seg_2_3_lutff_2_out_7010),
    .O(seg_2_3_local_g2_2_11575)
  );
  LocalMux t1753 (
    .I(seg_2_4_neigh_op_bot_2_7010),
    .O(seg_2_4_local_g0_2_11682)
  );
  LocalMux t1754 (
    .I(seg_2_2_neigh_op_top_3_7011),
    .O(seg_2_2_local_g0_3_11437)
  );
  LocalMux t1755 (
    .I(seg_2_4_neigh_op_bot_3_7011),
    .O(seg_2_4_local_g0_3_11683)
  );
  LocalMux t1756 (
    .I(seg_2_3_lutff_4_out_7012),
    .O(seg_2_3_local_g3_4_11585)
  );
  LocalMux t1757 (
    .I(seg_2_3_lutff_5_out_7013),
    .O(seg_2_3_local_g3_5_11586)
  );
  LocalMux t1758 (
    .I(seg_2_2_neigh_op_top_6_7014),
    .O(seg_2_2_local_g1_6_11448)
  );
  LocalMux t1759 (
    .I(seg_2_3_lutff_7_out_7015),
    .O(seg_2_3_local_g0_7_11564)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t176 (
    .carryinitin(),
    .carryinitout(t175)
  );
  LocalMux t1760 (
    .I(seg_6_4_sp4_h_r_45_15615),
    .O(seg_6_4_local_g2_5_26960)
  );
  Span4Mux_h3 t1761 (
    .I(seg_3_4_sp4_v_b_8_11421),
    .O(seg_6_4_sp4_h_r_45_15615)
  );
  LocalMux t1762 (
    .I(seg_6_4_sp4_h_r_47_15607),
    .O(seg_6_4_local_g2_7_26962)
  );
  Span4Mux_h3 t1763 (
    .I(seg_3_4_sp4_v_b_10_11423),
    .O(seg_6_4_sp4_h_r_47_15607)
  );
  LocalMux t1764 (
    .I(seg_2_4_lutff_0_out_7155),
    .O(seg_2_4_local_g2_0_11696)
  );
  LocalMux t1765 (
    .I(seg_1_3_neigh_op_tnr_1_7156),
    .O(seg_1_3_local_g2_1_7066)
  );
  LocalMux t1766 (
    .I(seg_1_4_neigh_op_rgt_1_7156),
    .O(seg_1_4_local_g2_1_7213)
  );
  LocalMux t1767 (
    .I(seg_1_4_neigh_op_rgt_2_7157),
    .O(seg_1_4_local_g2_2_7214)
  );
  LocalMux t1768 (
    .I(seg_2_4_lutff_2_out_7157),
    .O(seg_2_4_local_g3_2_11706)
  );
  LocalMux t1769 (
    .I(seg_2_3_neigh_op_top_3_7158),
    .O(seg_2_3_local_g0_3_11560)
  );
  LocalMux t1770 (
    .I(seg_2_4_lutff_4_out_7159),
    .O(seg_2_4_local_g1_4_11692)
  );
  LocalMux t1771 (
    .I(seg_2_3_neigh_op_top_5_7160),
    .O(seg_2_3_local_g1_5_11570)
  );
  LocalMux t1772 (
    .I(seg_3_4_neigh_op_lft_5_7160),
    .O(seg_3_4_local_g1_5_15524)
  );
  LocalMux t1773 (
    .I(seg_1_4_neigh_op_rgt_6_7161),
    .O(seg_1_4_local_g3_6_7226)
  );
  LocalMux t1774 (
    .I(seg_3_4_neigh_op_lft_6_7161),
    .O(seg_3_4_local_g1_6_15525)
  );
  LocalMux t1775 (
    .I(seg_3_4_neigh_op_lft_7_7162),
    .O(seg_3_4_local_g0_7_15518)
  );
  LocalMux t1776 (
    .I(seg_6_3_sp4_v_b_23_22916),
    .O(seg_6_3_local_g0_7_26844)
  );
  Span4Mux_v1 t1777 (
    .I(seg_6_4_sp4_h_l_47_11776),
    .O(seg_6_3_sp4_v_b_23_22916)
  );
  LocalMux t1778 (
    .I(seg_2_1_sp4_v_b_47_6891),
    .O(seg_2_1_local_g2_7_11294)
  );
  LocalMux t1779 (
    .I(seg_1_4_neigh_op_tnr_2_7304),
    .O(seg_1_4_local_g3_2_7222)
  );
  LocalMux t1780 (
    .I(seg_2_5_lutff_2_out_7304),
    .O(seg_2_5_local_g3_2_11829)
  );
  LocalMux t1781 (
    .I(seg_1_5_neigh_op_rgt_4_7306),
    .O(seg_1_5_local_g2_4_7363)
  );
  LocalMux t1782 (
    .I(seg_2_4_neigh_op_top_6_7308),
    .O(seg_2_4_local_g0_6_11686)
  );
  LocalMux t1783 (
    .I(seg_2_5_lutff_6_out_7308),
    .O(seg_2_5_local_g3_6_11833)
  );
  LocalMux t1784 (
    .I(seg_1_5_neigh_op_rgt_7_7309),
    .O(seg_1_5_local_g2_7_7366)
  );
  LocalMux t1785 (
    .I(seg_0_17_sp4_v_b_8_2930),
    .O(seg_0_17_local_g0_0_3580)
  );
  Span4Mux_v4 t1786 (
    .I(seg_0_13_sp4_v_b_8_2097),
    .O(seg_0_17_sp4_v_b_8_2930)
  );
  Span4Mux_v4 t1787 (
    .I(seg_0_9_sp4_v_b_8_1247),
    .O(seg_0_13_sp4_v_b_8_2097)
  );
  Span4Mux_v4 t1788 (
    .I(seg_0_5_sp4_h_r_8_1224),
    .O(seg_0_9_sp4_v_b_8_1247)
  );
  LocalMux t1789 (
    .I(seg_6_3_sp4_h_r_47_15484),
    .O(seg_6_3_local_g2_7_26860)
  );
  Span4Mux_h3 t1790 (
    .I(seg_3_3_sp4_v_t_40_11790),
    .O(seg_6_3_sp4_h_r_47_15484)
  );
  LocalMux t1791 (
    .I(seg_7_4_sp4_h_r_7_30307),
    .O(seg_7_4_local_g0_7_30211)
  );
  Span4Mux_h0 t1792 (
    .I(seg_7_4_sp4_h_l_42_15614),
    .O(seg_7_4_sp4_h_r_7_30307)
  );
  Span4Mux_h4 t1793 (
    .I(seg_3_4_sp4_v_t_39_11912),
    .O(seg_7_4_sp4_h_l_42_15614)
  );
  LocalMux t1794 (
    .I(seg_2_2_sp4_v_b_4_6858),
    .O(seg_2_2_local_g1_4_11446)
  );
  Span4Mux_v0 t1795 (
    .I(seg_2_2_sp4_v_t_36_7179),
    .O(seg_2_2_sp4_v_b_4_6858)
  );
  LocalMux t1796 (
    .I(seg_0_7_sp4_h_r_25_1610),
    .O(seg_0_7_local_g3_1_1485)
  );
  Span4Mux_h2 t1797 (
    .I(seg_2_7_sp4_v_b_8_7335),
    .O(seg_0_7_sp4_h_r_25_1610)
  );
  LocalMux t1798 (
    .I(seg_1_6_neigh_op_rgt_0_7449),
    .O(seg_1_6_local_g2_0_7506)
  );
  LocalMux t1799 (
    .I(seg_1_6_neigh_op_rgt_3_7452),
    .O(seg_1_6_local_g2_3_7509)
  );
  CascadeMux t18 (
    .I(net_7120),
    .O(net_7120_cascademuxed)
  );
  LocalMux t1800 (
    .I(seg_1_6_neigh_op_rgt_4_7453),
    .O(seg_1_6_local_g2_4_7510)
  );
  LocalMux t1801 (
    .I(seg_3_5_neigh_op_tnl_5_7454),
    .O(seg_3_5_local_g2_5_15655)
  );
  LocalMux t1802 (
    .I(seg_5_5_sp4_r_v_b_23_23167),
    .O(seg_5_5_local_g3_7_23327)
  );
  Span4Mux_v1 t1803 (
    .I(seg_6_6_sp4_h_l_47_12022),
    .O(seg_5_5_sp4_r_v_b_23_23167)
  );
  LocalMux t1804 (
    .I(seg_0_17_sp4_r_v_b_19_3353),
    .O(seg_0_17_local_g3_3_3607)
  );
  Span4Mux_v3 t1805 (
    .I(seg_1_14_sp4_v_b_3_2494),
    .O(seg_0_17_sp4_r_v_b_19_3353)
  );
  Span4Mux_v4 t1806 (
    .I(seg_1_10_sp4_v_b_3_1642),
    .O(seg_1_14_sp4_v_b_3_2494)
  );
  Span4Mux_v4 t1807 (
    .I(seg_1_6_sp4_h_r_9_7619),
    .O(seg_1_10_sp4_v_b_3_1642)
  );
  LocalMux t1808 (
    .I(seg_7_13_sp4_r_v_b_12_31171),
    .O(seg_7_13_local_g2_4_31331)
  );
  Span4Mux_v3 t1809 (
    .I(seg_8_10_sp4_v_b_1_30679),
    .O(seg_7_13_sp4_r_v_b_12_31171)
  );
  Span4Mux_v4 t1810 (
    .I(seg_8_6_sp4_h_l_36_19683),
    .O(seg_8_10_sp4_v_b_1_30679)
  );
  Span4Mux_h4 t1811 (
    .I(seg_4_6_sp4_h_l_47_1386),
    .O(seg_8_6_sp4_h_l_36_19683)
  );
  LocalMux t1812 (
    .I(seg_7_7_sp4_h_r_3_30672),
    .O(seg_7_7_local_g1_3_30584)
  );
  Span4Mux_h0 t1813 (
    .I(seg_7_7_sp4_h_l_37_15974),
    .O(seg_7_7_sp4_h_r_3_30672)
  );
  Span4Mux_h4 t1814 (
    .I(seg_3_7_sp4_v_b_0_11787),
    .O(seg_7_7_sp4_h_l_37_15974)
  );
  LocalMux t1815 (
    .I(seg_0_7_sp4_h_r_12_1596),
    .O(seg_0_7_local_g0_4_1464)
  );
  Span4Mux_h3 t1816 (
    .I(seg_3_7_sp4_v_b_8_11795),
    .O(seg_0_7_sp4_h_r_12_1596)
  );
  LocalMux t1817 (
    .I(seg_2_7_lutff_0_out_7596),
    .O(seg_2_7_local_g3_0_12073)
  );
  LocalMux t1818 (
    .I(seg_2_8_neigh_op_bot_3_7599),
    .O(seg_2_8_local_g0_3_12175)
  );
  LocalMux t1819 (
    .I(seg_2_8_neigh_op_bot_4_7600),
    .O(seg_2_8_local_g0_4_12176)
  );
  LocalMux t1820 (
    .I(seg_2_8_neigh_op_bot_6_7602),
    .O(seg_2_8_local_g1_6_12186)
  );
  LocalMux t1821 (
    .I(seg_2_8_neigh_op_bot_7_7603),
    .O(seg_2_8_local_g1_7_12187)
  );
  LocalMux t1822 (
    .I(seg_3_18_sp4_v_b_16_13266),
    .O(seg_3_18_local_g0_0_17233)
  );
  Span4Mux_v3 t1823 (
    .I(seg_3_15_sp4_v_b_9_12778),
    .O(seg_3_18_sp4_v_b_16_13266)
  );
  Span4Mux_v4 t1824 (
    .I(seg_3_11_sp4_v_b_6_12285),
    .O(seg_3_15_sp4_v_b_9_12778)
  );
  Span4Mux_v4 t1825 (
    .I(seg_3_7_sp4_v_b_3_11788),
    .O(seg_3_11_sp4_v_b_6_12285)
  );
  LocalMux t1826 (
    .I(seg_2_8_lutff_2_out_7745),
    .O(seg_2_8_local_g2_2_12190)
  );
  LocalMux t1827 (
    .I(seg_2_8_lutff_5_out_7748),
    .O(seg_2_8_local_g0_5_12177)
  );
  LocalMux t1828 (
    .I(seg_2_8_lutff_6_out_7749),
    .O(seg_2_8_local_g2_6_12194)
  );
  LocalMux t1829 (
    .I(seg_2_8_lutff_7_out_7750),
    .O(seg_2_8_local_g0_7_12179)
  );
  CascadeMux t183 (
    .I(net_16038),
    .O(net_16038_cascademuxed)
  );
  LocalMux t1830 (
    .I(seg_5_16_sp4_r_v_b_2_24389),
    .O(seg_5_16_local_g1_2_24659)
  );
  Span4Mux_v4 t1831 (
    .I(seg_6_12_sp4_v_b_6_23901),
    .O(seg_5_16_sp4_r_v_b_2_24389)
  );
  Span4Mux_v4 t1832 (
    .I(seg_6_8_sp4_h_l_43_12274),
    .O(seg_6_12_sp4_v_b_6_23901)
  );
  LocalMux t1833 (
    .I(seg_5_16_sp4_r_v_b_4_24391),
    .O(seg_5_16_local_g1_4_24661)
  );
  Span4Mux_v4 t1834 (
    .I(seg_6_12_sp4_v_b_1_23894),
    .O(seg_5_16_sp4_r_v_b_4_24391)
  );
  Span4Mux_v4 t1835 (
    .I(seg_6_8_sp4_h_l_45_12276),
    .O(seg_6_12_sp4_v_b_1_23894)
  );
  LocalMux t1836 (
    .I(seg_3_18_sp4_v_b_9_13147),
    .O(seg_3_18_local_g1_1_17242)
  );
  Span4Mux_v4 t1837 (
    .I(seg_3_14_sp4_v_b_9_12655),
    .O(seg_3_18_sp4_v_b_9_13147)
  );
  Span4Mux_v4 t1838 (
    .I(seg_3_10_sp4_v_b_9_12163),
    .O(seg_3_14_sp4_v_b_9_12655)
  );
  LocalMux t1839 (
    .I(seg_3_18_sp4_v_b_5_13143),
    .O(seg_3_18_local_g1_5_17246)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t184 (
    .carryinitin(net_19908),
    .carryinitout(net_19952)
  );
  Span4Mux_v4 t1840 (
    .I(seg_3_14_sp4_v_b_2_12650),
    .O(seg_3_18_sp4_v_b_5_13143)
  );
  Span4Mux_v4 t1841 (
    .I(seg_3_10_sp4_v_b_11_12165),
    .O(seg_3_14_sp4_v_b_2_12650)
  );
  LocalMux t1842 (
    .I(seg_2_9_lutff_0_out_7890),
    .O(seg_2_9_local_g0_0_12295)
  );
  LocalMux t1843 (
    .I(seg_3_8_neigh_op_tnl_1_7891),
    .O(seg_3_8_local_g2_1_16020)
  );
  LocalMux t1844 (
    .I(seg_3_9_neigh_op_lft_1_7891),
    .O(seg_3_9_local_g1_1_16135)
  );
  LocalMux t1845 (
    .I(seg_2_9_lutff_2_out_7892),
    .O(seg_2_9_local_g0_2_12297)
  );
  LocalMux t1846 (
    .I(seg_3_8_neigh_op_tnl_4_7894),
    .O(seg_3_8_local_g2_4_16023)
  );
  LocalMux t1847 (
    .I(seg_3_9_neigh_op_lft_4_7894),
    .O(seg_3_9_local_g1_4_16138)
  );
  LocalMux t1848 (
    .I(seg_3_9_neigh_op_lft_5_7895),
    .O(seg_3_9_local_g1_5_16139)
  );
  LocalMux t1849 (
    .I(seg_2_8_neigh_op_top_6_7896),
    .O(seg_2_8_local_g0_6_12178)
  );
  CascadeMux t185 (
    .I(net_16161),
    .O(net_16161_cascademuxed)
  );
  LocalMux t1850 (
    .I(seg_7_9_sp4_h_r_25_23883),
    .O(seg_7_9_local_g2_1_30836)
  );
  Span4Mux_h2 t1851 (
    .I(seg_5_9_sp4_h_l_36_8050),
    .O(seg_7_9_sp4_h_r_25_23883)
  );
  LocalMux t1852 (
    .I(seg_4_7_sp4_r_v_b_29_19698),
    .O(seg_4_7_local_g1_5_19724)
  );
  Span4Mux_v2 t1853 (
    .I(seg_5_9_sp4_h_l_46_8052),
    .O(seg_4_7_sp4_r_v_b_29_19698)
  );
  LocalMux t1854 (
    .I(seg_5_10_sp4_h_r_30_16351),
    .O(seg_5_10_local_g2_6_23933)
  );
  Span4Mux_h2 t1855 (
    .I(seg_3_10_sp4_v_b_0_12156),
    .O(seg_5_10_sp4_h_r_30_16351)
  );
  LocalMux t1856 (
    .I(seg_12_10_sp4_h_r_20_46371),
    .O(seg_12_10_local_g0_4_50101)
  );
  Span4Mux_h1 t1857 (
    .I(seg_11_10_sp4_h_l_44_31047),
    .O(seg_12_10_sp4_h_r_20_46371)
  );
  Span4Mux_h4 t1858 (
    .I(seg_7_10_sp4_h_l_43_16351),
    .O(seg_11_10_sp4_h_l_44_31047)
  );
  Span4Mux_h4 t1859 (
    .I(seg_3_10_sp4_v_b_0_12156),
    .O(seg_7_10_sp4_h_l_43_16351)
  );
  CascadeMux t186 (
    .I(net_16167),
    .O(net_16167_cascademuxed)
  );
  LocalMux t1860 (
    .I(seg_3_6_sp4_h_r_10_15853),
    .O(seg_3_6_local_g1_2_15767)
  );
  Span4Mux_h0 t1861 (
    .I(seg_3_6_sp4_v_t_47_12166),
    .O(seg_3_6_sp4_h_r_10_15853)
  );
  LocalMux t1862 (
    .I(seg_5_10_sp4_h_r_34_16345),
    .O(seg_5_10_local_g3_2_23937)
  );
  Span4Mux_h2 t1863 (
    .I(seg_3_10_sp4_v_b_10_12166),
    .O(seg_5_10_sp4_h_r_34_16345)
  );
  LocalMux t1864 (
    .I(seg_14_10_sp4_h_r_36_46361),
    .O(seg_14_10_local_g3_4_57786)
  );
  Span4Mux_h3 t1865 (
    .I(seg_11_10_sp4_h_l_36_31037),
    .O(seg_14_10_sp4_h_r_36_46361)
  );
  Span4Mux_h4 t1866 (
    .I(seg_7_10_sp4_h_l_47_16345),
    .O(seg_11_10_sp4_h_l_36_31037)
  );
  Span4Mux_h4 t1867 (
    .I(seg_3_10_sp4_v_b_10_12166),
    .O(seg_7_10_sp4_h_l_47_16345)
  );
  LocalMux t1868 (
    .I(seg_0_11_sp4_h_r_13_2449),
    .O(seg_0_11_local_g1_5_2327)
  );
  Span4Mux_h3 t1869 (
    .I(seg_3_11_sp4_v_b_7_12284),
    .O(seg_0_11_sp4_h_r_13_2449)
  );
  CascadeMux t187 (
    .I(net_16173),
    .O(net_16173_cascademuxed)
  );
  LocalMux t1870 (
    .I(seg_4_12_sp4_h_r_15_16593),
    .O(seg_4_12_local_g1_7_20341)
  );
  Span4Mux_h1 t1871 (
    .I(seg_3_12_sp4_v_b_2_12404),
    .O(seg_4_12_sp4_h_r_15_16593)
  );
  LocalMux t1872 (
    .I(seg_2_7_sp4_v_b_36_7767),
    .O(seg_2_7_local_g3_4_12077)
  );
  LocalMux t1873 (
    .I(seg_0_16_sp4_h_r_28_3525),
    .O(seg_0_16_local_g2_4_3394)
  );
  Span4Mux_h2 t1874 (
    .I(seg_2_16_sp4_v_b_11_8659),
    .O(seg_0_16_sp4_h_r_28_3525)
  );
  Span4Mux_v4 t1875 (
    .I(seg_2_12_sp4_v_b_11_8071),
    .O(seg_2_16_sp4_v_b_11_8659)
  );
  LocalMux t1876 (
    .I(seg_3_9_neigh_op_tnl_0_8037),
    .O(seg_3_9_local_g2_0_16142)
  );
  LocalMux t1877 (
    .I(seg_2_10_lutff_2_out_8039),
    .O(seg_2_10_local_g2_2_12436)
  );
  LocalMux t1878 (
    .I(seg_2_11_neigh_op_bot_4_8041),
    .O(seg_2_11_local_g1_4_12553)
  );
  LocalMux t1879 (
    .I(seg_3_9_neigh_op_tnl_6_8043),
    .O(seg_3_9_local_g3_6_16156)
  );
  CascadeMux t188 (
    .I(net_16179),
    .O(net_16179_cascademuxed)
  );
  LocalMux t1880 (
    .I(seg_3_9_neigh_op_tnl_7_8044),
    .O(seg_3_9_local_g2_7_16149)
  );
  LocalMux t1881 (
    .I(seg_3_18_sp4_v_b_0_13140),
    .O(seg_3_18_local_g1_0_17241)
  );
  Span4Mux_v4 t1882 (
    .I(seg_3_14_sp4_v_b_0_12648),
    .O(seg_3_18_sp4_v_b_0_13140)
  );
  Span4Mux_v4 t1883 (
    .I(seg_3_10_sp4_h_l_42_2248),
    .O(seg_3_14_sp4_v_b_0_12648)
  );
  LocalMux t1884 (
    .I(seg_3_12_sp4_v_b_13_12525),
    .O(seg_3_12_local_g0_5_16500)
  );
  LocalMux t1885 (
    .I(seg_1_10_neigh_op_tnr_1_8185),
    .O(seg_1_10_local_g2_1_8095)
  );
  LocalMux t1886 (
    .I(seg_1_10_neigh_op_tnr_2_8186),
    .O(seg_1_10_local_g3_2_8104)
  );
  LocalMux t1887 (
    .I(seg_1_11_neigh_op_rgt_3_8187),
    .O(seg_1_11_local_g3_3_8252)
  );
  LocalMux t1888 (
    .I(seg_3_11_neigh_op_lft_5_8189),
    .O(seg_3_11_local_g1_5_16385)
  );
  LocalMux t1889 (
    .I(seg_1_10_neigh_op_tnr_6_8190),
    .O(seg_1_10_local_g3_6_8108)
  );
  CascadeMux t189 (
    .I(net_16185),
    .O(net_16185_cascademuxed)
  );
  LocalMux t1890 (
    .I(seg_3_13_sp4_v_b_7_12530),
    .O(seg_3_13_local_g1_7_16633)
  );
  LocalMux t1891 (
    .I(seg_2_13_sp4_r_v_b_23_12658),
    .O(seg_2_13_local_g3_7_12818)
  );
  LocalMux t1892 (
    .I(seg_2_9_sp4_v_b_32_7923),
    .O(seg_2_9_local_g3_0_12319)
  );
  LocalMux t1893 (
    .I(seg_3_13_neigh_op_bnl_0_8331),
    .O(seg_3_13_local_g3_0_16642)
  );
  LocalMux t1894 (
    .I(seg_3_13_neigh_op_bnl_1_8332),
    .O(seg_3_13_local_g3_1_16643)
  );
  LocalMux t1895 (
    .I(seg_3_13_neigh_op_bnl_2_8333),
    .O(seg_3_13_local_g2_2_16636)
  );
  LocalMux t1896 (
    .I(seg_3_13_neigh_op_bnl_3_8334),
    .O(seg_3_13_local_g2_3_16637)
  );
  LocalMux t1897 (
    .I(seg_3_13_neigh_op_bnl_4_8335),
    .O(seg_3_13_local_g2_4_16638)
  );
  LocalMux t1898 (
    .I(seg_3_13_neigh_op_bnl_5_8336),
    .O(seg_3_13_local_g3_5_16647)
  );
  LocalMux t1899 (
    .I(seg_3_13_neigh_op_bnl_6_8337),
    .O(seg_3_13_local_g3_6_16648)
  );
  CascadeMux t19 (
    .I(net_7126),
    .O(net_7126_cascademuxed)
  );
  CascadeMux t190 (
    .I(net_16191),
    .O(net_16191_cascademuxed)
  );
  LocalMux t1900 (
    .I(seg_3_14_sp4_v_b_7_12653),
    .O(seg_3_14_local_g1_7_16756)
  );
  LocalMux t1901 (
    .I(seg_3_14_neigh_op_bnl_0_8478),
    .O(seg_3_14_local_g3_0_16765)
  );
  LocalMux t1902 (
    .I(seg_2_13_lutff_1_out_8479),
    .O(seg_2_13_local_g3_1_12812)
  );
  LocalMux t1903 (
    .I(seg_3_12_neigh_op_tnl_4_8482),
    .O(seg_3_12_local_g3_4_16523)
  );
  LocalMux t1904 (
    .I(seg_3_12_neigh_op_tnl_6_8484),
    .O(seg_3_12_local_g2_6_16517)
  );
  LocalMux t1905 (
    .I(seg_2_13_lutff_7_out_8485),
    .O(seg_2_13_local_g2_7_12810)
  );
  LocalMux t1906 (
    .I(seg_14_10_sp4_v_b_36_54034),
    .O(seg_14_10_local_g2_4_57778)
  );
  Span4Mux_v3 t1907 (
    .I(seg_14_13_sp4_h_l_36_42899),
    .O(seg_14_10_sp4_v_b_36_54034)
  );
  Span4Mux_h4 t1908 (
    .I(seg_10_13_sp4_h_l_36_27932),
    .O(seg_14_13_sp4_h_l_36_42899)
  );
  Span4Mux_h4 t1909 (
    .I(seg_6_13_sp4_h_l_47_12883),
    .O(seg_10_13_sp4_h_l_36_27932)
  );
  CascadeMux t191 (
    .I(net_16197),
    .O(net_16197_cascademuxed)
  );
  LocalMux t1910 (
    .I(seg_4_12_sp4_v_b_15_16358),
    .O(seg_4_12_local_g0_7_20333)
  );
  Span4Mux_v1 t1911 (
    .I(seg_4_13_sp4_h_l_39_2873),
    .O(seg_4_12_sp4_v_b_15_16358)
  );
  LocalMux t1912 (
    .I(seg_4_13_sp4_h_r_28_12887),
    .O(seg_4_13_local_g3_4_20477)
  );
  LocalMux t1913 (
    .I(seg_4_13_sp4_h_r_30_12889),
    .O(seg_4_13_local_g2_6_20471)
  );
  LocalMux t1914 (
    .I(seg_3_8_sp4_v_b_18_12038),
    .O(seg_3_8_local_g0_2_16005)
  );
  Span4Mux_v1 t1915 (
    .I(seg_3_9_sp4_v_t_46_12534),
    .O(seg_3_8_sp4_v_b_18_12038)
  );
  LocalMux t1916 (
    .I(seg_2_7_sp4_v_b_30_7627),
    .O(seg_2_7_local_g2_6_12071)
  );
  Span4Mux_v2 t1917 (
    .I(seg_2_9_sp4_v_t_47_8219),
    .O(seg_2_7_sp4_v_b_30_7627)
  );
  LocalMux t1918 (
    .I(seg_2_8_sp4_v_b_12_7620),
    .O(seg_2_8_local_g1_4_12184)
  );
  Span4Mux_v1 t1919 (
    .I(seg_2_9_sp4_v_t_47_8219),
    .O(seg_2_8_sp4_v_b_12_7620)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t192 (
    .carryinitin(net_20031),
    .carryinitout(net_20075)
  );
  LocalMux t1920 (
    .I(seg_2_10_sp4_h_r_1_12513),
    .O(seg_2_10_local_g0_1_12419)
  );
  Span4Mux_h0 t1921 (
    .I(seg_2_10_sp4_v_t_36_8355),
    .O(seg_2_10_sp4_h_r_1_12513)
  );
  LocalMux t1922 (
    .I(seg_4_14_sp4_h_r_34_13006),
    .O(seg_4_14_local_g3_2_20598)
  );
  LocalMux t1923 (
    .I(seg_7_14_sp4_h_r_25_24498),
    .O(seg_7_14_local_g3_1_31459)
  );
  Span4Mux_h2 t1924 (
    .I(seg_5_14_sp4_h_l_36_8785),
    .O(seg_7_14_sp4_h_r_25_24498)
  );
  LocalMux t1925 (
    .I(seg_7_13_sp4_v_b_20_27747),
    .O(seg_7_13_local_g0_4_31315)
  );
  Span4Mux_v1 t1926 (
    .I(seg_7_14_sp4_h_l_44_16846),
    .O(seg_7_13_sp4_v_b_20_27747)
  );
  Span4Mux_h4 t1927 (
    .I(seg_3_14_sp4_h_l_36_3092),
    .O(seg_7_14_sp4_h_l_44_16846)
  );
  LocalMux t1928 (
    .I(seg_3_10_sp4_v_b_27_12403),
    .O(seg_3_10_local_g2_3_16268)
  );
  Span4Mux_v2 t1929 (
    .I(seg_3_12_sp4_v_t_42_12899),
    .O(seg_3_10_sp4_v_b_27_12403)
  );
  CascadeMux t193 (
    .I(net_16296),
    .O(net_16296_cascademuxed)
  );
  LocalMux t1930 (
    .I(seg_5_12_sp4_h_r_35_16592),
    .O(seg_5_12_local_g3_3_24184)
  );
  Span4Mux_h2 t1931 (
    .I(seg_3_12_sp4_v_t_46_12903),
    .O(seg_5_12_sp4_h_r_35_16592)
  );
  LocalMux t1932 (
    .I(seg_3_10_sp4_h_r_19_12520),
    .O(seg_3_10_local_g1_3_16260)
  );
  Span4Mux_h1 t1933 (
    .I(seg_2_10_sp4_v_t_43_8362),
    .O(seg_3_10_sp4_h_r_19_12520)
  );
  LocalMux t1934 (
    .I(seg_2_9_sp4_v_b_21_7776),
    .O(seg_2_9_local_g1_5_12308)
  );
  Span4Mux_v1 t1935 (
    .I(seg_2_10_sp4_v_t_45_8364),
    .O(seg_2_9_sp4_v_b_21_7776)
  );
  LocalMux t1936 (
    .I(seg_2_14_neigh_op_top_1_8773),
    .O(seg_2_14_local_g1_1_12919)
  );
  LocalMux t1937 (
    .I(seg_2_14_neigh_op_top_2_8774),
    .O(seg_2_14_local_g1_2_12920)
  );
  LocalMux t1938 (
    .I(seg_2_14_neigh_op_top_3_8775),
    .O(seg_2_14_local_g0_3_12913)
  );
  LocalMux t1939 (
    .I(seg_2_15_lutff_4_out_8776),
    .O(seg_2_15_local_g0_4_13037)
  );
  CascadeMux t194 (
    .I(net_16320),
    .O(net_16320_cascademuxed)
  );
  LocalMux t1940 (
    .I(seg_3_15_neigh_op_lft_6_8778),
    .O(seg_3_15_local_g1_6_16878)
  );
  LocalMux t1941 (
    .I(seg_4_15_sp4_h_r_34_13129),
    .O(seg_4_15_local_g3_2_20721)
  );
  LocalMux t1942 (
    .I(seg_4_15_sp4_h_r_38_8936),
    .O(seg_4_15_local_g2_6_20717)
  );
  LocalMux t1943 (
    .I(seg_2_16_lutff_0_out_8919),
    .O(seg_2_16_local_g1_0_13164)
  );
  LocalMux t1944 (
    .I(seg_2_15_neigh_op_top_1_8920),
    .O(seg_2_15_local_g0_1_13034)
  );
  LocalMux t1945 (
    .I(seg_2_15_neigh_op_top_2_8921),
    .O(seg_2_15_local_g0_2_13035)
  );
  LocalMux t1946 (
    .I(seg_3_16_neigh_op_lft_3_8922),
    .O(seg_3_16_local_g1_3_16998)
  );
  LocalMux t1947 (
    .I(seg_3_15_neigh_op_tnl_4_8923),
    .O(seg_3_15_local_g2_4_16884)
  );
  LocalMux t1948 (
    .I(seg_3_15_neigh_op_tnl_5_8924),
    .O(seg_3_15_local_g3_5_16893)
  );
  LocalMux t1949 (
    .I(seg_2_15_neigh_op_top_6_8925),
    .O(seg_2_15_local_g0_6_13039)
  );
  CascadeMux t195 (
    .I(net_16326),
    .O(net_16326_cascademuxed)
  );
  LocalMux t1950 (
    .I(seg_2_15_neigh_op_top_7_8926),
    .O(seg_2_15_local_g0_7_13040)
  );
  LocalMux t1951 (
    .I(seg_2_16_neigh_op_top_2_9068),
    .O(seg_2_16_local_g1_2_13166)
  );
  LocalMux t1952 (
    .I(seg_3_16_neigh_op_tnl_5_9071),
    .O(seg_3_16_local_g3_5_17016)
  );
  LocalMux t1953 (
    .I(seg_2_16_neigh_op_top_7_9073),
    .O(seg_2_16_local_g0_7_13163)
  );
  LocalMux t1954 (
    .I(seg_3_17_neigh_op_tnl_0_9213),
    .O(seg_3_17_local_g2_0_17126)
  );
  LocalMux t1955 (
    .I(seg_3_17_neigh_op_tnl_1_9214),
    .O(seg_3_17_local_g2_1_17127)
  );
  LocalMux t1956 (
    .I(seg_2_17_neigh_op_top_4_9217),
    .O(seg_2_17_local_g1_4_13291)
  );
  LocalMux t1957 (
    .I(seg_3_17_neigh_op_tnl_6_9219),
    .O(seg_3_17_local_g2_6_17132)
  );
  LocalMux t1958 (
    .I(seg_3_17_neigh_op_tnl_7_9220),
    .O(seg_3_17_local_g2_7_17133)
  );
  LocalMux t1959 (
    .I(seg_3_19_neigh_op_lft_0_9360),
    .O(seg_3_19_local_g1_0_17364)
  );
  CascadeMux t196 (
    .I(net_16419),
    .O(net_16419_cascademuxed)
  );
  LocalMux t1960 (
    .I(seg_2_18_neigh_op_top_1_9361),
    .O(seg_2_18_local_g0_1_13403)
  );
  LocalMux t1961 (
    .I(seg_3_18_neigh_op_tnl_4_9364),
    .O(seg_3_18_local_g2_4_17253)
  );
  LocalMux t1962 (
    .I(seg_2_18_neigh_op_top_5_9365),
    .O(seg_2_18_local_g0_5_13407)
  );
  LocalMux t1963 (
    .I(seg_2_19_lutff_6_out_9366),
    .O(seg_2_19_local_g0_6_13531)
  );
  LocalMux t1964 (
    .I(seg_2_18_neigh_op_top_7_9367),
    .O(seg_2_18_local_g0_7_13409)
  );
  LocalMux t1965 (
    .I(seg_2_16_sp4_v_b_43_9097),
    .O(seg_2_16_local_g3_3_13183)
  );
  LocalMux t1966 (
    .I(seg_3_19_neigh_op_tnl_1_9508),
    .O(seg_3_19_local_g2_1_17373)
  );
  LocalMux t1967 (
    .I(seg_2_19_neigh_op_top_3_9510),
    .O(seg_2_19_local_g0_3_13528)
  );
  LocalMux t1968 (
    .I(seg_2_19_neigh_op_top_4_9511),
    .O(seg_2_19_local_g1_4_13537)
  );
  LocalMux t1969 (
    .I(seg_2_19_neigh_op_top_5_9512),
    .O(seg_2_19_local_g1_5_13538)
  );
  CascadeMux t197 (
    .I(net_16425),
    .O(net_16425_cascademuxed)
  );
  LocalMux t1970 (
    .I(seg_2_19_neigh_op_top_7_9514),
    .O(seg_2_19_local_g1_7_13540)
  );
  LocalMux t1971 (
    .I(seg_2_20_neigh_op_top_4_9658),
    .O(seg_2_20_local_g0_4_13652)
  );
  LocalMux t1972 (
    .I(seg_2_17_sp4_h_r_7_13382),
    .O(seg_2_17_local_g1_7_13294)
  );
  Span4Mux_h0 t1973 (
    .I(seg_2_17_sp4_v_t_39_9387),
    .O(seg_2_17_sp4_h_r_7_13382)
  );
  LocalMux t1974 (
    .I(seg_2_21_neigh_op_top_0_9801),
    .O(seg_2_21_local_g1_0_13779)
  );
  LocalMux t1975 (
    .I(seg_2_21_neigh_op_top_5_9806),
    .O(seg_2_21_local_g0_5_13776)
  );
  LocalMux t1976 (
    .I(seg_3_22_neigh_op_tnl_4_9952),
    .O(seg_3_22_local_g2_4_17745)
  );
  LocalMux t1977 (
    .I(seg_3_1_lutff_0_out_11229),
    .O(seg_3_1_local_g2_0_15118)
  );
  LocalMux t1978 (
    .I(seg_3_1_lutff_1_out_11230),
    .O(seg_3_1_local_g0_1_15103)
  );
  LocalMux t1979 (
    .I(seg_4_2_neigh_op_bnl_1_11230),
    .O(seg_4_2_local_g2_1_19113)
  );
  CascadeMux t198 (
    .I(net_16431),
    .O(net_16431_cascademuxed)
  );
  LocalMux t1980 (
    .I(seg_4_1_neigh_op_lft_2_11231),
    .O(seg_4_1_local_g1_2_18943)
  );
  LocalMux t1981 (
    .I(seg_4_2_neigh_op_bnl_2_11231),
    .O(seg_4_2_local_g2_2_19114)
  );
  LocalMux t1982 (
    .I(seg_4_1_neigh_op_lft_3_11232),
    .O(seg_4_1_local_g0_3_18936)
  );
  LocalMux t1983 (
    .I(seg_4_2_neigh_op_bnl_3_11232),
    .O(seg_4_2_local_g3_3_19123)
  );
  LocalMux t1984 (
    .I(seg_2_1_neigh_op_rgt_6_11235),
    .O(seg_2_1_local_g2_6_11293)
  );
  LocalMux t1985 (
    .I(seg_2_2_neigh_op_bnr_6_11235),
    .O(seg_2_2_local_g0_6_11440)
  );
  LocalMux t1986 (
    .I(seg_4_1_neigh_op_lft_7_11236),
    .O(seg_4_1_local_g1_7_18948)
  );
  LocalMux t1987 (
    .I(seg_4_2_neigh_op_bnl_7_11236),
    .O(seg_4_2_local_g2_7_19119)
  );
  LocalMux t1988 (
    .I(seg_6_4_sp4_v_b_19_23040),
    .O(seg_6_4_local_g1_3_26950)
  );
  Span4Mux_v3 t1989 (
    .I(seg_6_1_sp4_h_l_36_11370),
    .O(seg_6_4_sp4_v_b_19_23040)
  );
  CascadeMux t199 (
    .I(net_16443),
    .O(net_16443_cascademuxed)
  );
  LocalMux t1990 (
    .I(seg_6_4_sp4_v_b_14_23035),
    .O(seg_6_4_local_g0_6_26945)
  );
  Span4Mux_v3 t1991 (
    .I(seg_6_1_sp4_h_l_38_11374),
    .O(seg_6_4_sp4_v_b_14_23035)
  );
  LocalMux t1992 (
    .I(seg_6_4_sp4_v_b_18_23039),
    .O(seg_6_4_local_g1_2_26949)
  );
  Span4Mux_v3 t1993 (
    .I(seg_6_1_sp4_h_l_42_11378),
    .O(seg_6_4_sp4_v_b_18_23039)
  );
  LocalMux t1994 (
    .I(seg_6_4_sp4_v_b_20_23041),
    .O(seg_6_4_local_g0_4_26943)
  );
  Span4Mux_v3 t1995 (
    .I(seg_6_1_sp4_h_l_44_11380),
    .O(seg_6_4_sp4_v_b_20_23041)
  );
  LocalMux t1996 (
    .I(seg_1_1_sp4_h_r_20_250),
    .O(seg_1_1_local_g1_4_6727)
  );
  LocalMux t1997 (
    .I(seg_6_4_sp4_r_v_b_22_26831),
    .O(seg_6_4_local_g3_6_26969)
  );
  Span4Mux_v3 t1998 (
    .I(seg_7_1_sp4_h_l_43_15208),
    .O(seg_6_4_sp4_r_v_b_22_26831)
  );
  LocalMux t1999 (
    .I(seg_1_3_sp4_h_r_23_743),
    .O(seg_1_3_local_g0_7_7056)
  );
  CascadeMux t20 (
    .I(net_7231),
    .O(net_7231_cascademuxed)
  );
  CascadeMux t200 (
    .I(net_16530),
    .O(net_16530_cascademuxed)
  );
  Span4Mux_h3 t2000 (
    .I(seg_4_3_sp4_v_b_5_15234),
    .O(seg_1_3_sp4_h_r_23_743)
  );
  LocalMux t2001 (
    .I(seg_5_3_sp4_h_r_22_19316),
    .O(seg_5_3_local_g0_6_23056)
  );
  Span4Mux_h1 t2002 (
    .I(seg_4_3_sp4_v_b_5_15234),
    .O(seg_5_3_sp4_h_r_22_19316)
  );
  LocalMux t2003 (
    .I(seg_3_2_lutff_0_out_11357),
    .O(seg_3_2_local_g3_0_15289)
  );
  LocalMux t2004 (
    .I(seg_3_2_lutff_1_out_11358),
    .O(seg_3_2_local_g1_1_15274)
  );
  LocalMux t2005 (
    .I(seg_3_2_lutff_2_out_11359),
    .O(seg_3_2_local_g3_2_15291)
  );
  LocalMux t2006 (
    .I(seg_4_2_neigh_op_lft_2_11359),
    .O(seg_4_2_local_g0_2_19098)
  );
  LocalMux t2007 (
    .I(seg_3_2_lutff_3_out_11360),
    .O(seg_3_2_local_g2_3_15284)
  );
  LocalMux t2008 (
    .I(seg_3_2_lutff_4_out_11361),
    .O(seg_3_2_local_g0_4_15269)
  );
  LocalMux t2009 (
    .I(seg_4_2_neigh_op_lft_4_11361),
    .O(seg_4_2_local_g1_4_19108)
  );
  CascadeMux t201 (
    .I(net_16536),
    .O(net_16536_cascademuxed)
  );
  LocalMux t2010 (
    .I(seg_3_2_lutff_5_out_11362),
    .O(seg_3_2_local_g3_5_15294)
  );
  LocalMux t2011 (
    .I(seg_3_2_lutff_6_out_11363),
    .O(seg_3_2_local_g3_6_15295)
  );
  LocalMux t2012 (
    .I(seg_3_3_neigh_op_bot_6_11363),
    .O(seg_3_3_local_g0_6_15394)
  );
  LocalMux t2013 (
    .I(seg_4_3_neigh_op_bnl_6_11363),
    .O(seg_4_3_local_g2_6_19241)
  );
  LocalMux t2014 (
    .I(seg_3_2_lutff_7_out_11364),
    .O(seg_3_2_local_g3_7_15296)
  );
  LocalMux t2015 (
    .I(seg_4_2_neigh_op_lft_7_11364),
    .O(seg_4_2_local_g0_7_19103)
  );
  LocalMux t2016 (
    .I(seg_6_4_sp4_r_v_b_28_26928),
    .O(seg_6_4_local_g1_4_26951)
  );
  Span4Mux_v2 t2017 (
    .I(seg_7_2_sp4_h_l_41_15365),
    .O(seg_6_4_sp4_r_v_b_28_26928)
  );
  LocalMux t2018 (
    .I(seg_6_4_sp4_r_v_b_32_26932),
    .O(seg_6_4_local_g2_0_26955)
  );
  Span4Mux_v2 t2019 (
    .I(seg_7_2_sp4_h_l_45_15369),
    .O(seg_6_4_sp4_r_v_b_32_26932)
  );
  CascadeMux t202 (
    .I(net_16542),
    .O(net_16542_cascademuxed)
  );
  LocalMux t2020 (
    .I(seg_6_3_sp4_h_r_30_19321),
    .O(seg_6_3_local_g3_6_26867)
  );
  Span4Mux_h2 t2021 (
    .I(seg_4_3_sp4_v_b_0_15229),
    .O(seg_6_3_sp4_h_r_30_19321)
  );
  LocalMux t2022 (
    .I(seg_6_4_sp4_h_r_25_19437),
    .O(seg_6_4_local_g3_1_26964)
  );
  Span4Mux_h2 t2023 (
    .I(seg_4_4_sp4_v_b_7_15249),
    .O(seg_6_4_sp4_h_r_25_19437)
  );
  LocalMux t2024 (
    .I(seg_3_2_neigh_op_top_0_11516),
    .O(seg_3_2_local_g1_0_15273)
  );
  LocalMux t2025 (
    .I(seg_3_3_lutff_1_out_11517),
    .O(seg_3_3_local_g1_1_15397)
  );
  LocalMux t2026 (
    .I(seg_3_3_lutff_2_out_11518),
    .O(seg_3_3_local_g1_2_15398)
  );
  LocalMux t2027 (
    .I(seg_4_3_neigh_op_lft_2_11518),
    .O(seg_4_3_local_g0_2_19221)
  );
  LocalMux t2028 (
    .I(seg_3_3_lutff_3_out_11519),
    .O(seg_3_3_local_g1_3_15399)
  );
  LocalMux t2029 (
    .I(seg_4_3_neigh_op_lft_3_11519),
    .O(seg_4_3_local_g0_3_19222)
  );
  CascadeMux t203 (
    .I(net_16548),
    .O(net_16548_cascademuxed)
  );
  LocalMux t2030 (
    .I(seg_3_3_lutff_4_out_11520),
    .O(seg_3_3_local_g3_4_15416)
  );
  LocalMux t2031 (
    .I(seg_4_3_neigh_op_lft_4_11520),
    .O(seg_4_3_local_g0_4_19223)
  );
  LocalMux t2032 (
    .I(seg_3_3_lutff_5_out_11521),
    .O(seg_3_3_local_g2_5_15409)
  );
  LocalMux t2033 (
    .I(seg_3_3_lutff_6_out_11522),
    .O(seg_3_3_local_g1_6_15402)
  );
  LocalMux t2034 (
    .I(seg_3_3_lutff_7_out_11523),
    .O(seg_3_3_local_g0_7_15395)
  );
  LocalMux t2035 (
    .I(seg_6_3_sp4_h_r_41_15488),
    .O(seg_6_3_local_g3_1_26862)
  );
  LocalMux t2036 (
    .I(seg_6_3_sp4_h_r_43_15490),
    .O(seg_6_3_local_g2_3_26856)
  );
  LocalMux t2037 (
    .I(seg_6_4_sp4_r_v_b_29_26927),
    .O(seg_6_4_local_g0_5_26944)
  );
  Span4Mux_v2 t2038 (
    .I(seg_7_6_sp4_h_l_40_15858),
    .O(seg_6_4_sp4_r_v_b_29_26927)
  );
  Span4Mux_h4 t2039 (
    .I(seg_3_6_sp4_v_b_5_11667),
    .O(seg_7_6_sp4_h_l_40_15858)
  );
  CascadeMux t204 (
    .I(net_16554),
    .O(net_16554_cascademuxed)
  );
  LocalMux t2040 (
    .I(seg_3_4_lutff_0_out_11639),
    .O(seg_3_4_local_g1_0_15519)
  );
  LocalMux t2041 (
    .I(seg_3_5_neigh_op_bot_0_11639),
    .O(seg_3_5_local_g1_0_15642)
  );
  LocalMux t2042 (
    .I(seg_4_5_neigh_op_bnl_0_11639),
    .O(seg_4_5_local_g2_0_19481)
  );
  LocalMux t2043 (
    .I(seg_3_3_neigh_op_top_2_11641),
    .O(seg_3_3_local_g0_2_15390)
  );
  LocalMux t2044 (
    .I(seg_4_3_neigh_op_tnl_2_11641),
    .O(seg_4_3_local_g2_2_19237)
  );
  LocalMux t2045 (
    .I(seg_4_3_neigh_op_tnl_2_11641),
    .O(seg_4_3_local_g3_2_19245)
  );
  LocalMux t2046 (
    .I(seg_4_4_neigh_op_lft_2_11641),
    .O(seg_4_4_local_g1_2_19352)
  );
  LocalMux t2047 (
    .I(seg_2_4_neigh_op_rgt_3_11642),
    .O(seg_2_4_local_g3_3_11707)
  );
  LocalMux t2048 (
    .I(seg_3_4_lutff_3_out_11642),
    .O(seg_3_4_local_g0_3_15514)
  );
  LocalMux t2049 (
    .I(seg_2_4_neigh_op_rgt_4_11643),
    .O(seg_2_4_local_g3_4_11708)
  );
  CascadeMux t205 (
    .I(net_16560),
    .O(net_16560_cascademuxed)
  );
  LocalMux t2050 (
    .I(seg_3_4_lutff_4_out_11643),
    .O(seg_3_4_local_g1_4_15523)
  );
  LocalMux t2051 (
    .I(seg_3_4_lutff_5_out_11644),
    .O(seg_3_4_local_g0_5_15516)
  );
  LocalMux t2052 (
    .I(seg_2_4_neigh_op_rgt_6_11645),
    .O(seg_2_4_local_g2_6_11702)
  );
  LocalMux t2053 (
    .I(seg_2_3_neigh_op_tnr_7_11646),
    .O(seg_2_3_local_g3_7_11588)
  );
  LocalMux t2054 (
    .I(seg_6_3_sp4_v_b_12_22904),
    .O(seg_6_3_local_g0_4_26841)
  );
  Span4Mux_v1 t2055 (
    .I(seg_6_4_sp4_h_l_36_11775),
    .O(seg_6_3_sp4_v_b_12_22904)
  );
  LocalMux t2056 (
    .I(seg_4_7_sp4_v_b_17_15745),
    .O(seg_4_7_local_g0_1_19712)
  );
  Span4Mux_v3 t2057 (
    .I(seg_4_4_sp4_v_b_1_15242),
    .O(seg_4_7_sp4_v_b_17_15745)
  );
  LocalMux t2058 (
    .I(seg_4_7_sp4_v_b_17_15745),
    .O(seg_4_7_local_g1_1_19720)
  );
  LocalMux t2059 (
    .I(seg_3_2_sp4_r_v_b_29_15247),
    .O(seg_3_2_local_g0_5_15270)
  );
  CascadeMux t206 (
    .I(net_16566),
    .O(net_16566_cascademuxed)
  );
  LocalMux t2060 (
    .I(seg_3_2_sp4_r_v_b_34_15254),
    .O(seg_3_2_local_g2_2_15283)
  );
  Span4Mux_v2 t2061 (
    .I(seg_4_4_sp4_h_l_47_970),
    .O(seg_3_2_sp4_r_v_b_34_15254)
  );
  Span4Mux_h0 t2062 (
    .I(seg_4_4_sp4_v_b_5_15247),
    .O(seg_4_4_sp4_h_l_47_970)
  );
  LocalMux t2063 (
    .I(seg_4_1_sp4_v_b_40_15247),
    .O(seg_4_1_local_g2_0_18949)
  );
  LocalMux t2064 (
    .I(seg_3_1_sp4_h_r_2_15204),
    .O(seg_3_1_local_g0_2_15104)
  );
  Span4Mux_h0 t2065 (
    .I(seg_3_1_sp4_v_t_44_11548),
    .O(seg_3_1_sp4_h_r_2_15204)
  );
  LocalMux t2066 (
    .I(seg_2_2_sp4_h_r_47_530),
    .O(seg_2_2_local_g3_7_11465)
  );
  Span4Mux_h1 t2067 (
    .I(seg_3_2_sp4_v_t_41_11668),
    .O(seg_2_2_sp4_h_r_47_530)
  );
  LocalMux t2068 (
    .I(seg_3_6_sp4_v_b_8_11672),
    .O(seg_3_6_local_g1_0_15765)
  );
  LocalMux t2069 (
    .I(seg_3_1_sp4_v_b_41_11417),
    .O(seg_3_1_local_g2_1_15119)
  );
  LocalMux t2070 (
    .I(seg_3_1_sp4_v_b_41_11417),
    .O(seg_3_1_local_g3_1_15127)
  );
  LocalMux t2071 (
    .I(seg_2_4_neigh_op_tnr_0_11762),
    .O(seg_2_4_local_g3_0_11704)
  );
  LocalMux t2072 (
    .I(seg_2_5_neigh_op_rgt_0_11762),
    .O(seg_2_5_local_g2_0_11819)
  );
  LocalMux t2073 (
    .I(seg_3_4_neigh_op_top_0_11762),
    .O(seg_3_4_local_g0_0_15511)
  );
  LocalMux t2074 (
    .I(seg_4_4_neigh_op_tnl_2_11764),
    .O(seg_4_4_local_g2_2_19360)
  );
  LocalMux t2075 (
    .I(seg_2_5_neigh_op_rgt_4_11766),
    .O(seg_2_5_local_g3_4_11831)
  );
  LocalMux t2076 (
    .I(seg_2_5_neigh_op_rgt_6_11768),
    .O(seg_2_5_local_g2_6_11825)
  );
  LocalMux t2077 (
    .I(seg_9_5_sp4_h_r_1_38084),
    .O(seg_9_5_local_g1_1_37998)
  );
  Span4Mux_h0 t2078 (
    .I(seg_9_5_sp4_h_l_40_23397),
    .O(seg_9_5_sp4_h_r_1_38084)
  );
  Span4Mux_h4 t2079 (
    .I(seg_5_5_sp4_h_l_39_7465),
    .O(seg_9_5_sp4_h_l_40_23397)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t208 (
    .carryinitin(),
    .carryinitout(t207)
  );
  LocalMux t2080 (
    .I(seg_1_5_sp4_h_r_6_7469),
    .O(seg_1_5_local_g0_6_7349)
  );
  LocalMux t2081 (
    .I(seg_1_3_sp4_v_b_25_562),
    .O(seg_1_3_local_g3_1_7074)
  );
  Span4Mux_v2 t2082 (
    .I(seg_1_5_sp4_h_r_8_7471),
    .O(seg_1_3_sp4_v_b_25_562)
  );
  LocalMux t2083 (
    .I(seg_1_5_sp4_h_r_8_7471),
    .O(seg_1_5_local_g0_0_7343)
  );
  LocalMux t2084 (
    .I(seg_1_5_sp4_h_r_10_7463),
    .O(seg_1_5_local_g1_2_7353)
  );
  LocalMux t2085 (
    .I(seg_6_3_sp4_h_r_26_19317),
    .O(seg_6_3_local_g2_2_26855)
  );
  Span4Mux_h2 t2086 (
    .I(seg_4_3_sp4_v_t_44_15625),
    .O(seg_6_3_sp4_h_r_26_19317)
  );
  LocalMux t2087 (
    .I(seg_2_1_sp4_r_v_b_0_11381),
    .O(seg_2_1_local_g1_0_11279)
  );
  Span4Mux_v1 t2088 (
    .I(seg_3_1_sp4_v_t_37_11541),
    .O(seg_2_1_sp4_r_v_b_0_11381)
  );
  LocalMux t2089 (
    .I(seg_4_6_neigh_op_lft_0_11885),
    .O(seg_4_6_local_g1_0_19596)
  );
  LocalMux t2090 (
    .I(seg_3_6_lutff_1_out_11886),
    .O(seg_3_6_local_g2_1_15774)
  );
  LocalMux t2091 (
    .I(seg_4_7_neigh_op_bnl_5_11890),
    .O(seg_4_7_local_g3_5_19740)
  );
  LocalMux t2092 (
    .I(seg_4_7_neigh_op_bnl_7_11892),
    .O(seg_4_7_local_g2_7_19734)
  );
  LocalMux t2093 (
    .I(seg_5_17_sp4_r_v_b_12_24632),
    .O(seg_5_17_local_g2_4_24792)
  );
  Span4Mux_v3 t2094 (
    .I(seg_6_14_sp4_v_b_1_24140),
    .O(seg_5_17_sp4_r_v_b_12_24632)
  );
  Span4Mux_v4 t2095 (
    .I(seg_6_10_sp4_v_b_1_23648),
    .O(seg_6_14_sp4_v_b_1_24140)
  );
  Span4Mux_v4 t2096 (
    .I(seg_6_6_sp4_h_l_36_12021),
    .O(seg_6_10_sp4_v_b_1_23648)
  );
  LocalMux t2097 (
    .I(seg_15_6_sp4_v_b_2_57006),
    .O(seg_15_6_local_g0_2_61098)
  );
  Span4Mux_v0 t2098 (
    .I(seg_15_6_sp4_h_l_45_45878),
    .O(seg_15_6_sp4_v_b_2_57006)
  );
  Span4Mux_h4 t2099 (
    .I(seg_11_6_sp4_h_l_45_30554),
    .O(seg_15_6_sp4_h_l_45_45878)
  );
  CascadeMux t21 (
    .I(net_7261),
    .O(net_7261_cascademuxed)
  );
  Span4Mux_h4 t2100 (
    .I(seg_7_6_sp4_h_l_45_15861),
    .O(seg_11_6_sp4_h_l_45_30554)
  );
  LocalMux t2101 (
    .I(seg_5_7_sp4_h_r_29_15981),
    .O(seg_5_7_local_g3_5_23571)
  );
  Span4Mux_h2 t2102 (
    .I(seg_3_7_sp4_v_b_11_11796),
    .O(seg_5_7_sp4_h_r_29_15981)
  );
  LocalMux t2103 (
    .I(seg_2_6_neigh_op_tnr_1_12009),
    .O(seg_2_6_local_g2_1_11943)
  );
  LocalMux t2104 (
    .I(seg_2_6_neigh_op_tnr_4_12012),
    .O(seg_2_6_local_g3_4_11954)
  );
  LocalMux t2105 (
    .I(seg_2_6_neigh_op_tnr_6_12014),
    .O(seg_2_6_local_g3_6_11956)
  );
  LocalMux t2106 (
    .I(seg_2_6_neigh_op_tnr_7_12015),
    .O(seg_2_6_local_g3_7_11957)
  );
  LocalMux t2107 (
    .I(seg_1_8_sp4_v_b_39_1852),
    .O(seg_1_8_local_g3_7_7815)
  );
  Span4Mux_v1 t2108 (
    .I(seg_1_7_sp4_h_r_2_7759),
    .O(seg_1_8_sp4_v_b_39_1852)
  );
  LocalMux t2109 (
    .I(seg_5_12_sp4_h_r_24_16589),
    .O(seg_5_12_local_g2_0_24173)
  );
  Span4Mux_h2 t2110 (
    .I(seg_3_12_sp4_v_b_0_12402),
    .O(seg_5_12_sp4_h_r_24_16589)
  );
  Span4Mux_v4 t2111 (
    .I(seg_3_8_sp4_v_b_9_11917),
    .O(seg_3_12_sp4_v_b_0_12402)
  );
  LocalMux t2112 (
    .I(seg_1_8_sp4_h_r_28_1810),
    .O(seg_1_8_local_g3_4_7812)
  );
  Span4Mux_h2 t2113 (
    .I(seg_3_8_sp4_v_b_11_11919),
    .O(seg_1_8_sp4_h_r_28_1810)
  );
  LocalMux t2114 (
    .I(seg_4_8_neigh_op_lft_4_12135),
    .O(seg_4_8_local_g0_4_19838)
  );
  LocalMux t2115 (
    .I(seg_5_16_sp4_r_v_b_5_24390),
    .O(seg_5_16_local_g1_5_24662)
  );
  Span4Mux_v4 t2116 (
    .I(seg_6_12_sp4_v_b_2_23897),
    .O(seg_5_16_sp4_r_v_b_5_24390)
  );
  Span4Mux_v4 t2117 (
    .I(seg_6_8_sp4_h_l_44_12277),
    .O(seg_6_12_sp4_v_b_2_23897)
  );
  LocalMux t2118 (
    .I(seg_3_18_sp4_v_b_4_13144),
    .O(seg_3_18_local_g0_4_17237)
  );
  Span4Mux_v4 t2119 (
    .I(seg_3_14_sp4_v_b_8_12656),
    .O(seg_3_18_sp4_v_b_4_13144)
  );
  Span4Mux_v4 t2120 (
    .I(seg_3_10_sp4_v_b_8_12164),
    .O(seg_3_14_sp4_v_b_8_12656)
  );
  LocalMux t2121 (
    .I(seg_3_18_sp4_v_b_23_13273),
    .O(seg_3_18_local_g1_7_17248)
  );
  Span4Mux_v3 t2122 (
    .I(seg_3_15_sp4_v_b_7_12776),
    .O(seg_3_18_sp4_v_b_23_13273)
  );
  Span4Mux_v4 t2123 (
    .I(seg_3_11_sp4_v_b_11_12288),
    .O(seg_3_15_sp4_v_b_7_12776)
  );
  LocalMux t2124 (
    .I(seg_4_8_neigh_op_tnl_1_12255),
    .O(seg_4_8_local_g3_1_19859)
  );
  LocalMux t2125 (
    .I(seg_4_8_neigh_op_tnl_2_12256),
    .O(seg_4_8_local_g2_2_19852)
  );
  LocalMux t2126 (
    .I(seg_4_8_neigh_op_tnl_3_12257),
    .O(seg_4_8_local_g3_3_19861)
  );
  LocalMux t2127 (
    .I(seg_4_8_neigh_op_tnl_4_12258),
    .O(seg_4_8_local_g2_4_19854)
  );
  LocalMux t2128 (
    .I(seg_4_8_neigh_op_tnl_5_12259),
    .O(seg_4_8_local_g3_5_19863)
  );
  LocalMux t2129 (
    .I(seg_4_8_neigh_op_tnl_6_12260),
    .O(seg_4_8_local_g2_6_19856)
  );
  LocalMux t2130 (
    .I(seg_4_8_neigh_op_tnl_7_12261),
    .O(seg_4_8_local_g3_7_19865)
  );
  LocalMux t2131 (
    .I(seg_4_9_neigh_op_lft_7_12261),
    .O(seg_4_9_local_g1_7_19972)
  );
  LocalMux t2132 (
    .I(seg_4_10_neigh_op_bnl_7_12261),
    .O(seg_4_10_local_g3_7_20111)
  );
  LocalMux t2133 (
    .I(seg_3_9_neigh_op_top_0_12377),
    .O(seg_3_9_local_g1_0_16134)
  );
  LocalMux t2134 (
    .I(seg_3_9_neigh_op_top_1_12378),
    .O(seg_3_9_local_g0_1_16127)
  );
  LocalMux t2135 (
    .I(seg_3_9_neigh_op_top_3_12380),
    .O(seg_3_9_local_g0_3_16129)
  );
  LocalMux t2136 (
    .I(seg_3_9_neigh_op_top_4_12381),
    .O(seg_3_9_local_g0_4_16130)
  );
  LocalMux t2137 (
    .I(seg_3_10_lutff_5_out_12382),
    .O(seg_3_10_local_g3_5_16278)
  );
  LocalMux t2138 (
    .I(seg_3_9_neigh_op_top_7_12384),
    .O(seg_3_9_local_g1_7_16141)
  );
  LocalMux t2139 (
    .I(seg_11_7_sp4_v_b_42_42178),
    .O(seg_11_7_local_g3_2_45923)
  );
  Span4Mux_v3 t2140 (
    .I(seg_11_10_sp4_h_l_42_31045),
    .O(seg_11_7_sp4_v_b_42_42178)
  );
  Span4Mux_h4 t2141 (
    .I(seg_7_10_sp4_h_l_41_16349),
    .O(seg_11_10_sp4_h_l_42_31045)
  );
  LocalMux t2142 (
    .I(seg_14_10_sp4_h_r_47_46362),
    .O(seg_14_10_local_g2_7_57781)
  );
  Span4Mux_h3 t2143 (
    .I(seg_11_10_sp4_h_l_42_31045),
    .O(seg_14_10_sp4_h_r_47_46362)
  );
  LocalMux t2144 (
    .I(seg_7_4_sp4_h_r_45_19446),
    .O(seg_7_4_local_g2_5_30225)
  );
  Span4Mux_h3 t2145 (
    .I(seg_4_4_sp4_v_t_45_15749),
    .O(seg_7_4_sp4_h_r_45_19446)
  );
  Span4Mux_v4 t2146 (
    .I(seg_4_8_sp4_v_t_40_16236),
    .O(seg_4_4_sp4_v_t_45_15749)
  );
  LocalMux t2147 (
    .I(seg_3_6_sp4_h_r_9_15862),
    .O(seg_3_6_local_g1_1_15766)
  );
  Span4Mux_h0 t2148 (
    .I(seg_3_6_sp4_v_t_41_12160),
    .O(seg_3_6_sp4_h_r_9_15862)
  );
  LocalMux t2149 (
    .I(seg_4_6_sp4_h_r_20_15862),
    .O(seg_4_6_local_g0_4_19592)
  );
  CascadeMux t215 (
    .I(net_16653),
    .O(net_16653_cascademuxed)
  );
  Span4Mux_h1 t2150 (
    .I(seg_3_6_sp4_v_t_41_12160),
    .O(seg_4_6_sp4_h_r_20_15862)
  );
  LocalMux t2151 (
    .I(seg_5_6_sp4_h_r_33_15862),
    .O(seg_5_6_local_g2_1_23436)
  );
  Span4Mux_h2 t2152 (
    .I(seg_3_6_sp4_v_t_41_12160),
    .O(seg_5_6_sp4_h_r_33_15862)
  );
  LocalMux t2153 (
    .I(seg_3_11_lutff_2_out_12502),
    .O(seg_3_11_local_g2_2_16390)
  );
  LocalMux t2154 (
    .I(seg_3_10_neigh_op_top_4_12504),
    .O(seg_3_10_local_g0_4_16253)
  );
  LocalMux t2155 (
    .I(seg_3_12_neigh_op_bot_7_12507),
    .O(seg_3_12_local_g1_7_16510)
  );
  LocalMux t2156 (
    .I(seg_0_6_sp4_v_b_21_810),
    .O(seg_0_6_local_g0_5_1259)
  );
  Span4Mux_v1 t2157 (
    .I(seg_0_7_sp4_v_t_37_1653),
    .O(seg_0_6_sp4_v_b_21_810)
  );
  Span4Mux_v4 t2158 (
    .I(seg_0_11_sp4_h_r_7_2489),
    .O(seg_0_7_sp4_v_t_37_1653)
  );
  LocalMux t2159 (
    .I(seg_0_6_sp4_v_b_16_805),
    .O(seg_0_6_local_g1_0_1262)
  );
  CascadeMux t216 (
    .I(net_16659),
    .O(net_16659_cascademuxed)
  );
  Span4Mux_v1 t2160 (
    .I(seg_0_7_sp4_v_t_44_1660),
    .O(seg_0_6_sp4_v_b_16_805)
  );
  Span4Mux_v4 t2161 (
    .I(seg_0_11_sp4_h_r_9_2491),
    .O(seg_0_7_sp4_v_t_44_1660)
  );
  LocalMux t2162 (
    .I(seg_0_6_sp4_v_b_19_808),
    .O(seg_0_6_local_g0_3_1257)
  );
  Span4Mux_v1 t2163 (
    .I(seg_0_7_sp4_h_r_1_1593),
    .O(seg_0_6_sp4_v_b_19_808)
  );
  Span4Mux_h4 t2164 (
    .I(seg_4_7_sp4_v_t_36_16109),
    .O(seg_0_7_sp4_h_r_1_1593)
  );
  LocalMux t2165 (
    .I(seg_0_24_sp4_v_b_23_4673),
    .O(seg_0_24_local_g0_7_5122)
  );
  Span4Mux_v3 t2166 (
    .I(seg_0_21_sp4_h_r_4_4636),
    .O(seg_0_24_sp4_v_b_23_4673)
  );
  Span4Mux_h4 t2167 (
    .I(seg_4_21_sp4_v_b_11_17349),
    .O(seg_0_21_sp4_h_r_4_4636)
  );
  Span4Mux_v4 t2168 (
    .I(seg_4_17_sp4_v_b_3_16849),
    .O(seg_4_21_sp4_v_b_11_17349)
  );
  Span4Mux_v4 t2169 (
    .I(seg_4_13_sp4_v_b_3_16357),
    .O(seg_4_17_sp4_v_b_3_16849)
  );
  CascadeMux t217 (
    .I(net_16665),
    .O(net_16665_cascademuxed)
  );
  LocalMux t2170 (
    .I(seg_0_24_sp4_v_b_13_4663),
    .O(seg_0_24_local_g0_5_5120)
  );
  Span4Mux_v3 t2171 (
    .I(seg_0_21_sp4_v_b_0_3773),
    .O(seg_0_24_sp4_v_b_13_4663)
  );
  Span4Mux_v4 t2172 (
    .I(seg_0_17_sp4_h_r_6_3756),
    .O(seg_0_21_sp4_v_b_0_3773)
  );
  Span4Mux_h4 t2173 (
    .I(seg_4_17_sp4_v_b_1_16847),
    .O(seg_0_17_sp4_h_r_6_3756)
  );
  Span4Mux_v4 t2174 (
    .I(seg_4_13_sp4_v_b_5_16359),
    .O(seg_4_17_sp4_v_b_1_16847)
  );
  LocalMux t2175 (
    .I(seg_0_6_sp4_v_b_14_803),
    .O(seg_0_6_local_g1_6_1268)
  );
  Span4Mux_v1 t2176 (
    .I(seg_0_7_sp4_h_r_3_1615),
    .O(seg_0_6_sp4_v_b_14_803)
  );
  Span4Mux_h4 t2177 (
    .I(seg_4_7_sp4_v_t_38_16111),
    .O(seg_0_7_sp4_h_r_3_1615)
  );
  LocalMux t2178 (
    .I(seg_0_24_sp4_v_b_16_4666),
    .O(seg_0_24_local_g1_0_5123)
  );
  Span4Mux_v3 t2179 (
    .I(seg_0_21_sp4_v_b_2_3775),
    .O(seg_0_24_sp4_v_b_16_4666)
  );
  CascadeMux t218 (
    .I(net_16671),
    .O(net_16671_cascademuxed)
  );
  Span4Mux_v4 t2180 (
    .I(seg_0_17_sp4_h_r_2_3724),
    .O(seg_0_21_sp4_v_b_2_3775)
  );
  Span4Mux_h4 t2181 (
    .I(seg_4_17_sp4_v_b_9_16855),
    .O(seg_0_17_sp4_h_r_2_3724)
  );
  Span4Mux_v4 t2182 (
    .I(seg_4_13_sp4_v_b_9_16363),
    .O(seg_4_17_sp4_v_b_9_16855)
  );
  LocalMux t2183 (
    .I(seg_0_6_sp4_v_b_18_807),
    .O(seg_0_6_local_g1_2_1264)
  );
  Span4Mux_v1 t2184 (
    .I(seg_0_7_sp4_h_r_7_1637),
    .O(seg_0_6_sp4_v_b_18_807)
  );
  Span4Mux_h4 t2185 (
    .I(seg_4_7_sp4_v_t_42_16115),
    .O(seg_0_7_sp4_h_r_7_1637)
  );
  LocalMux t2186 (
    .I(seg_0_24_sp4_h_r_18_5255),
    .O(seg_0_24_local_g1_2_5125)
  );
  Span4Mux_h3 t2187 (
    .I(seg_3_24_sp4_v_b_2_13880),
    .O(seg_0_24_sp4_h_r_18_5255)
  );
  Span4Mux_v4 t2188 (
    .I(seg_3_20_sp4_v_b_6_13392),
    .O(seg_3_24_sp4_v_b_2_13880)
  );
  Span4Mux_v4 t2189 (
    .I(seg_3_16_sp4_v_b_10_12904),
    .O(seg_3_20_sp4_v_b_6_13392)
  );
  CascadeMux t219 (
    .I(net_16677),
    .O(net_16677_cascademuxed)
  );
  Span4Mux_v4 t2190 (
    .I(seg_3_12_sp4_v_b_7_12407),
    .O(seg_3_16_sp4_v_b_10_12904)
  );
  LocalMux t2191 (
    .I(seg_0_24_sp4_h_r_12_5249),
    .O(seg_0_24_local_g1_4_5127)
  );
  Span4Mux_h3 t2192 (
    .I(seg_3_24_sp4_v_b_8_13886),
    .O(seg_0_24_sp4_h_r_12_5249)
  );
  Span4Mux_v4 t2193 (
    .I(seg_3_20_sp4_v_b_5_13389),
    .O(seg_3_24_sp4_v_b_8_13886)
  );
  Span4Mux_v4 t2194 (
    .I(seg_3_16_sp4_v_b_2_12896),
    .O(seg_3_20_sp4_v_b_5_13389)
  );
  Span4Mux_v4 t2195 (
    .I(seg_3_12_sp4_v_b_11_12411),
    .O(seg_3_16_sp4_v_b_2_12896)
  );
  LocalMux t2196 (
    .I(seg_2_11_neigh_op_tnr_1_12624),
    .O(seg_2_11_local_g3_1_12566)
  );
  LocalMux t2197 (
    .I(seg_2_11_neigh_op_tnr_2_12625),
    .O(seg_2_11_local_g2_2_12559)
  );
  LocalMux t2198 (
    .I(seg_2_11_neigh_op_tnr_3_12626),
    .O(seg_2_11_local_g3_3_12568)
  );
  LocalMux t2199 (
    .I(seg_2_11_neigh_op_tnr_4_12627),
    .O(seg_2_11_local_g3_4_12569)
  );
  CascadeMux t22 (
    .I(net_7273),
    .O(net_7273_cascademuxed)
  );
  CascadeMux t220 (
    .I(net_16683),
    .O(net_16683_cascademuxed)
  );
  LocalMux t2200 (
    .I(seg_2_11_neigh_op_tnr_5_12628),
    .O(seg_2_11_local_g3_5_12570)
  );
  LocalMux t2201 (
    .I(seg_2_11_neigh_op_tnr_6_12629),
    .O(seg_2_11_local_g2_6_12563)
  );
  LocalMux t2202 (
    .I(seg_2_11_neigh_op_tnr_7_12630),
    .O(seg_2_11_local_g2_7_12564)
  );
  LocalMux t2203 (
    .I(seg_2_12_neigh_op_rgt_7_12630),
    .O(seg_2_12_local_g3_7_12695)
  );
  LocalMux t2204 (
    .I(seg_2_13_neigh_op_bnr_7_12630),
    .O(seg_2_13_local_g1_7_12802)
  );
  LocalMux t2205 (
    .I(seg_2_14_neigh_op_bnr_7_12753),
    .O(seg_2_14_local_g1_7_12925)
  );
  LocalMux t2206 (
    .I(seg_5_13_sp4_h_r_34_16714),
    .O(seg_5_13_local_g3_2_24306)
  );
  LocalMux t2207 (
    .I(seg_8_13_sp4_h_r_28_27937),
    .O(seg_8_13_local_g3_4_35170)
  );
  Span4Mux_h2 t2208 (
    .I(seg_6_13_sp4_h_l_36_12882),
    .O(seg_8_13_sp4_h_r_28_27937)
  );
  LocalMux t2209 (
    .I(seg_5_13_sp4_h_r_26_16716),
    .O(seg_5_13_local_g2_2_24298)
  );
  CascadeMux t221 (
    .I(net_16689),
    .O(net_16689_cascademuxed)
  );
  LocalMux t2210 (
    .I(seg_5_13_sp4_h_r_44_12892),
    .O(seg_5_13_local_g2_4_24300)
  );
  LocalMux t2211 (
    .I(seg_5_13_sp4_h_r_46_12884),
    .O(seg_5_13_local_g3_6_24310)
  );
  LocalMux t2212 (
    .I(seg_5_13_sp4_h_r_32_16722),
    .O(seg_5_13_local_g2_0_24296)
  );
  LocalMux t2213 (
    .I(seg_2_14_neigh_op_rgt_0_12869),
    .O(seg_2_14_local_g3_0_12934)
  );
  LocalMux t2214 (
    .I(seg_2_14_neigh_op_rgt_1_12870),
    .O(seg_2_14_local_g3_1_12935)
  );
  LocalMux t2215 (
    .I(seg_3_14_lutff_2_out_12871),
    .O(seg_3_14_local_g3_2_16767)
  );
  LocalMux t2216 (
    .I(seg_2_13_neigh_op_tnr_5_12874),
    .O(seg_2_13_local_g3_5_12816)
  );
  LocalMux t2217 (
    .I(seg_3_13_neigh_op_top_5_12874),
    .O(seg_3_13_local_g0_5_16623)
  );
  LocalMux t2218 (
    .I(seg_3_12_sp4_r_v_b_39_16604),
    .O(seg_3_12_local_g2_7_16518)
  );
  LocalMux t2219 (
    .I(seg_3_12_sp4_v_b_36_12770),
    .O(seg_3_12_local_g2_4_16515)
  );
  CascadeMux t222 (
    .I(net_16695),
    .O(net_16695_cascademuxed)
  );
  LocalMux t2220 (
    .I(seg_3_10_sp4_v_b_32_12410),
    .O(seg_3_10_local_g3_0_16273)
  );
  Span4Mux_v2 t2221 (
    .I(seg_3_12_sp4_v_t_37_12894),
    .O(seg_3_10_sp4_v_b_32_12410)
  );
  LocalMux t2222 (
    .I(seg_3_9_sp4_v_b_15_12158),
    .O(seg_3_9_local_g0_7_16133)
  );
  Span4Mux_v1 t2223 (
    .I(seg_3_10_sp4_v_t_43_12654),
    .O(seg_3_9_sp4_v_b_15_12158)
  );
  LocalMux t2224 (
    .I(seg_3_14_neigh_op_top_7_12999),
    .O(seg_3_14_local_g0_7_16748)
  );
  LocalMux t2225 (
    .I(seg_3_13_sp4_r_v_b_37_16725),
    .O(seg_3_13_local_g2_5_16639)
  );
  LocalMux t2226 (
    .I(seg_3_13_sp4_r_v_b_43_16731),
    .O(seg_3_13_local_g3_3_16645)
  );
  LocalMux t2227 (
    .I(seg_3_13_sp4_r_v_b_31_16607),
    .O(seg_3_13_local_g0_7_16625)
  );
  LocalMux t2228 (
    .I(seg_3_13_sp4_v_b_34_12781),
    .O(seg_3_13_local_g3_2_16644)
  );
  LocalMux t2229 (
    .I(seg_3_13_sp4_v_b_38_12895),
    .O(seg_3_13_local_g2_6_16640)
  );
  CascadeMux t223 (
    .I(net_16776),
    .O(net_16776_cascademuxed)
  );
  LocalMux t2230 (
    .I(seg_3_13_sp4_v_b_28_12775),
    .O(seg_3_13_local_g3_4_16646)
  );
  LocalMux t2231 (
    .I(seg_3_13_sp4_v_b_32_12779),
    .O(seg_3_13_local_g2_0_16634)
  );
  LocalMux t2232 (
    .I(seg_3_15_neigh_op_top_0_13115),
    .O(seg_3_15_local_g0_0_16864)
  );
  LocalMux t2233 (
    .I(seg_3_15_neigh_op_top_1_13116),
    .O(seg_3_15_local_g1_1_16873)
  );
  LocalMux t2234 (
    .I(seg_3_15_neigh_op_top_2_13117),
    .O(seg_3_15_local_g0_2_16866)
  );
  LocalMux t2235 (
    .I(seg_3_15_neigh_op_top_4_13119),
    .O(seg_3_15_local_g0_4_16868)
  );
  LocalMux t2236 (
    .I(seg_3_15_neigh_op_top_5_13120),
    .O(seg_3_15_local_g0_5_16869)
  );
  LocalMux t2237 (
    .I(seg_2_16_neigh_op_rgt_7_13122),
    .O(seg_2_16_local_g3_7_13187)
  );
  LocalMux t2238 (
    .I(seg_3_9_sp4_h_r_6_16228),
    .O(seg_3_9_local_g0_6_16132)
  );
  Span4Mux_h0 t2239 (
    .I(seg_3_9_sp4_v_t_36_12524),
    .O(seg_3_9_sp4_h_r_6_16228)
  );
  CascadeMux t224 (
    .I(net_16782),
    .O(net_16782_cascademuxed)
  );
  Span4Mux_v4 t2240 (
    .I(seg_3_13_sp4_v_t_36_13016),
    .O(seg_3_9_sp4_v_t_36_12524)
  );
  LocalMux t2241 (
    .I(seg_3_14_sp4_v_b_28_12898),
    .O(seg_3_14_local_g2_4_16761)
  );
  LocalMux t2242 (
    .I(seg_3_9_sp4_v_b_43_12408),
    .O(seg_3_9_local_g3_3_16153)
  );
  Span4Mux_v3 t2243 (
    .I(seg_3_12_sp4_v_t_43_12900),
    .O(seg_3_9_sp4_v_b_43_12408)
  );
  LocalMux t2244 (
    .I(seg_3_16_neigh_op_top_2_13240),
    .O(seg_3_16_local_g0_2_16989)
  );
  LocalMux t2245 (
    .I(seg_3_16_neigh_op_top_3_13241),
    .O(seg_3_16_local_g0_3_16990)
  );
  LocalMux t2246 (
    .I(seg_3_16_neigh_op_top_4_13242),
    .O(seg_3_16_local_g1_4_16999)
  );
  LocalMux t2247 (
    .I(seg_3_16_neigh_op_top_5_13243),
    .O(seg_3_16_local_g0_5_16992)
  );
  LocalMux t2248 (
    .I(seg_3_16_neigh_op_top_6_13244),
    .O(seg_3_16_local_g1_6_17001)
  );
  LocalMux t2249 (
    .I(seg_3_11_sp4_v_b_32_12533),
    .O(seg_3_11_local_g2_0_16388)
  );
  CascadeMux t225 (
    .I(net_16794),
    .O(net_16794_cascademuxed)
  );
  Span4Mux_v2 t2250 (
    .I(seg_3_13_sp4_v_t_37_13017),
    .O(seg_3_11_sp4_v_b_32_12533)
  );
  LocalMux t2251 (
    .I(seg_3_15_sp4_v_b_38_13141),
    .O(seg_3_15_local_g2_6_16886)
  );
  LocalMux t2252 (
    .I(seg_4_6_sp4_h_r_7_19691),
    .O(seg_4_6_local_g1_7_19603)
  );
  Span4Mux_h0 t2253 (
    .I(seg_4_6_sp4_v_t_42_15992),
    .O(seg_4_6_sp4_h_r_7_19691)
  );
  Span4Mux_v4 t2254 (
    .I(seg_4_10_sp4_v_t_41_16483),
    .O(seg_4_6_sp4_v_t_42_15992)
  );
  Span4Mux_v4 t2255 (
    .I(seg_4_14_sp4_v_t_36_16970),
    .O(seg_4_10_sp4_v_t_41_16483)
  );
  LocalMux t2256 (
    .I(seg_4_6_sp4_h_r_3_19687),
    .O(seg_4_6_local_g1_3_19599)
  );
  Span4Mux_h0 t2257 (
    .I(seg_4_6_sp4_v_t_38_15988),
    .O(seg_4_6_sp4_h_r_3_19687)
  );
  Span4Mux_v4 t2258 (
    .I(seg_4_10_sp4_v_t_42_16484),
    .O(seg_4_6_sp4_v_t_38_15988)
  );
  Span4Mux_v4 t2259 (
    .I(seg_4_14_sp4_v_t_46_16980),
    .O(seg_4_10_sp4_v_t_42_16484)
  );
  CascadeMux t226 (
    .I(net_16812),
    .O(net_16812_cascademuxed)
  );
  LocalMux t2260 (
    .I(seg_4_5_sp4_v_b_35_15627),
    .O(seg_4_5_local_g3_3_19492)
  );
  Span4Mux_v2 t2261 (
    .I(seg_4_7_sp4_v_t_46_16119),
    .O(seg_4_5_sp4_v_b_35_15627)
  );
  Span4Mux_v4 t2262 (
    .I(seg_4_11_sp4_v_t_45_16610),
    .O(seg_4_7_sp4_v_t_46_16119)
  );
  Span4Mux_v4 t2263 (
    .I(seg_4_15_sp4_v_t_37_17094),
    .O(seg_4_11_sp4_v_t_45_16610)
  );
  LocalMux t2264 (
    .I(seg_3_12_sp4_v_b_46_12780),
    .O(seg_3_12_local_g3_6_16525)
  );
  Span4Mux_v3 t2265 (
    .I(seg_3_15_sp4_v_t_38_13264),
    .O(seg_3_12_sp4_v_b_46_12780)
  );
  LocalMux t2266 (
    .I(seg_3_12_sp4_v_b_35_12657),
    .O(seg_3_12_local_g2_3_16514)
  );
  Span4Mux_v2 t2267 (
    .I(seg_3_14_sp4_v_t_45_13148),
    .O(seg_3_12_sp4_v_b_35_12657)
  );
  LocalMux t2268 (
    .I(seg_3_18_neigh_op_top_5_13489),
    .O(seg_3_18_local_g0_5_17238)
  );
  LocalMux t2269 (
    .I(seg_3_17_sp4_r_v_b_29_17097),
    .O(seg_3_17_local_g0_5_17115)
  );
  CascadeMux t227 (
    .I(net_16899),
    .O(net_16899_cascademuxed)
  );
  LocalMux t2270 (
    .I(seg_3_14_sp4_v_b_29_12897),
    .O(seg_3_14_local_g2_5_16762)
  );
  Span4Mux_v2 t2271 (
    .I(seg_3_16_sp4_v_t_39_13388),
    .O(seg_3_14_sp4_v_b_29_12897)
  );
  LocalMux t2272 (
    .I(seg_3_17_sp4_h_r_3_17209),
    .O(seg_3_17_local_g1_3_17121)
  );
  Span4Mux_h0 t2273 (
    .I(seg_3_17_sp4_v_t_47_13519),
    .O(seg_3_17_sp4_h_r_3_17209)
  );
  LocalMux t2274 (
    .I(seg_3_17_sp4_v_b_12_13139),
    .O(seg_3_17_local_g0_4_17114)
  );
  Span4Mux_v1 t2275 (
    .I(seg_3_18_sp4_v_t_36_13631),
    .O(seg_3_17_sp4_v_b_12_13139)
  );
  LocalMux t2276 (
    .I(seg_3_21_neigh_op_top_3_13856),
    .O(seg_3_21_local_g1_3_17613)
  );
  LocalMux t2277 (
    .I(seg_3_1_neigh_op_rgt_0_15060),
    .O(seg_3_1_local_g3_0_15126)
  );
  LocalMux t2278 (
    .I(seg_4_1_lutff_2_out_15062),
    .O(seg_4_1_local_g2_2_18951)
  );
  LocalMux t2279 (
    .I(seg_3_1_neigh_op_rgt_3_15063),
    .O(seg_3_1_local_g2_3_15121)
  );
  CascadeMux t228 (
    .I(net_16905),
    .O(net_16905_cascademuxed)
  );
  LocalMux t2280 (
    .I(seg_3_2_neigh_op_bnr_3_15063),
    .O(seg_3_2_local_g0_3_15268)
  );
  LocalMux t2281 (
    .I(seg_4_1_lutff_4_out_15064),
    .O(seg_4_1_local_g1_4_18945)
  );
  LocalMux t2282 (
    .I(seg_3_1_neigh_op_rgt_5_15065),
    .O(seg_3_1_local_g3_5_15131)
  );
  LocalMux t2283 (
    .I(seg_4_1_lutff_5_out_15065),
    .O(seg_4_1_local_g1_5_18946)
  );
  LocalMux t2284 (
    .I(seg_3_1_neigh_op_rgt_6_15066),
    .O(seg_3_1_local_g3_6_15132)
  );
  LocalMux t2285 (
    .I(seg_3_1_neigh_op_rgt_7_15067),
    .O(seg_3_1_local_g3_7_15133)
  );
  LocalMux t2286 (
    .I(seg_4_3_sp4_r_v_b_15_19076),
    .O(seg_4_3_local_g2_7_19242)
  );
  LocalMux t2287 (
    .I(seg_4_4_sp4_r_v_b_4_19079),
    .O(seg_4_4_local_g1_4_19354)
  );
  LocalMux t2288 (
    .I(seg_3_4_sp4_h_r_30_7322),
    .O(seg_3_4_local_g2_6_15533)
  );
  Span4Mux_h2 t2289 (
    .I(seg_5_4_sp4_v_b_6_19081),
    .O(seg_3_4_sp4_h_r_30_7322)
  );
  CascadeMux t229 (
    .I(net_16911),
    .O(net_16911_cascademuxed)
  );
  LocalMux t2290 (
    .I(seg_3_3_sp4_r_v_b_14_15244),
    .O(seg_3_3_local_g2_6_15410)
  );
  LocalMux t2291 (
    .I(seg_3_2_neigh_op_rgt_1_15189),
    .O(seg_3_2_local_g2_1_15282)
  );
  LocalMux t2292 (
    .I(seg_4_1_neigh_op_top_2_15190),
    .O(seg_4_1_local_g0_2_18935)
  );
  LocalMux t2293 (
    .I(seg_4_1_neigh_op_top_3_15191),
    .O(seg_4_1_local_g1_3_18944)
  );
  LocalMux t2294 (
    .I(seg_3_2_neigh_op_rgt_4_15192),
    .O(seg_3_2_local_g2_4_15285)
  );
  LocalMux t2295 (
    .I(seg_3_2_neigh_op_rgt_5_15193),
    .O(seg_3_2_local_g2_5_15286)
  );
  LocalMux t2296 (
    .I(seg_3_1_neigh_op_tnr_6_15194),
    .O(seg_3_1_local_g2_6_15124)
  );
  LocalMux t2297 (
    .I(seg_4_1_neigh_op_top_7_15195),
    .O(seg_4_1_local_g0_7_18940)
  );
  LocalMux t2298 (
    .I(seg_3_3_neigh_op_rgt_0_15347),
    .O(seg_3_3_local_g3_0_15412)
  );
  LocalMux t2299 (
    .I(seg_4_3_lutff_1_out_15348),
    .O(seg_4_3_local_g2_1_19236)
  );
  CascadeMux t23 (
    .I(net_7384),
    .O(net_7384_cascademuxed)
  );
  CascadeMux t230 (
    .I(net_16917),
    .O(net_16917_cascademuxed)
  );
  LocalMux t2300 (
    .I(seg_3_3_neigh_op_rgt_2_15349),
    .O(seg_3_3_local_g2_2_15406)
  );
  LocalMux t2301 (
    .I(seg_3_3_neigh_op_rgt_3_15350),
    .O(seg_3_3_local_g3_3_15415)
  );
  LocalMux t2302 (
    .I(seg_3_3_neigh_op_rgt_4_15351),
    .O(seg_3_3_local_g2_4_15408)
  );
  LocalMux t2303 (
    .I(seg_4_3_lutff_5_out_15352),
    .O(seg_4_3_local_g0_5_19224)
  );
  LocalMux t2304 (
    .I(seg_4_3_lutff_5_out_15352),
    .O(seg_4_3_local_g1_5_19232)
  );
  LocalMux t2305 (
    .I(seg_4_2_neigh_op_top_6_15353),
    .O(seg_4_2_local_g0_6_19102)
  );
  LocalMux t2306 (
    .I(seg_4_4_neigh_op_bot_6_15353),
    .O(seg_4_4_local_g1_6_19356)
  );
  LocalMux t2307 (
    .I(seg_4_3_lutff_7_out_15354),
    .O(seg_4_3_local_g3_7_19250)
  );
  LocalMux t2308 (
    .I(seg_6_3_sp4_h_r_14_23149),
    .O(seg_6_3_local_g0_6_26843)
  );
  Span4Mux_h1 t2309 (
    .I(seg_5_3_sp4_h_l_42_7176),
    .O(seg_6_3_sp4_h_r_14_23149)
  );
  CascadeMux t231 (
    .I(net_16923),
    .O(net_16923_cascademuxed)
  );
  LocalMux t2310 (
    .I(seg_3_3_neigh_op_tnr_0_15470),
    .O(seg_3_3_local_g2_0_15404)
  );
  LocalMux t2311 (
    .I(seg_3_4_neigh_op_rgt_0_15470),
    .O(seg_3_4_local_g2_0_15527)
  );
  LocalMux t2312 (
    .I(seg_4_4_lutff_0_out_15470),
    .O(seg_4_4_local_g1_0_19350)
  );
  LocalMux t2313 (
    .I(seg_3_3_neigh_op_tnr_3_15473),
    .O(seg_3_3_local_g2_3_15407)
  );
  LocalMux t2314 (
    .I(seg_3_4_neigh_op_rgt_3_15473),
    .O(seg_3_4_local_g2_3_15530)
  );
  LocalMux t2315 (
    .I(seg_4_3_neigh_op_top_3_15473),
    .O(seg_4_3_local_g1_3_19230)
  );
  LocalMux t2316 (
    .I(seg_4_4_lutff_3_out_15473),
    .O(seg_4_4_local_g1_3_19353)
  );
  LocalMux t2317 (
    .I(seg_4_4_lutff_3_out_15473),
    .O(seg_4_4_local_g2_3_19361)
  );
  LocalMux t2318 (
    .I(seg_4_4_lutff_4_out_15474),
    .O(seg_4_4_local_g2_4_19362)
  );
  LocalMux t2319 (
    .I(seg_4_3_neigh_op_top_6_15476),
    .O(seg_4_3_local_g0_6_19225)
  );
  CascadeMux t232 (
    .I(net_16929),
    .O(net_16929_cascademuxed)
  );
  LocalMux t2320 (
    .I(seg_7_3_sp4_r_v_b_15_29938),
    .O(seg_7_3_local_g2_7_30104)
  );
  Span4Mux_v1 t2321 (
    .I(seg_8_4_sp4_h_l_39_19440),
    .O(seg_7_3_sp4_r_v_b_15_29938)
  );
  LocalMux t2322 (
    .I(seg_8_4_sp4_h_r_29_27020),
    .O(seg_8_4_local_g2_5_34056)
  );
  Span4Mux_h2 t2323 (
    .I(seg_6_4_sp4_h_l_39_11778),
    .O(seg_8_4_sp4_h_r_29_27020)
  );
  LocalMux t2324 (
    .I(seg_7_3_sp4_r_v_b_23_29947),
    .O(seg_7_3_local_g3_7_30112)
  );
  Span4Mux_v1 t2325 (
    .I(seg_8_4_sp4_h_l_41_19442),
    .O(seg_7_3_sp4_r_v_b_23_29947)
  );
  LocalMux t2326 (
    .I(seg_5_1_sp4_v_b_42_19080),
    .O(seg_5_1_local_g3_2_22790)
  );
  LocalMux t2327 (
    .I(seg_3_2_sp4_r_v_b_24_15243),
    .O(seg_3_2_local_g0_0_15265)
  );
  LocalMux t2328 (
    .I(seg_4_1_sp4_v_b_37_15243),
    .O(seg_4_1_local_g2_5_18954)
  );
  LocalMux t2329 (
    .I(seg_4_1_sp4_v_b_43_15250),
    .O(seg_4_1_local_g2_3_18952)
  );
  CascadeMux t233 (
    .I(net_16935),
    .O(net_16935_cascademuxed)
  );
  LocalMux t2330 (
    .I(seg_4_2_sp4_v_b_30_15250),
    .O(seg_4_2_local_g2_6_19118)
  );
  LocalMux t2331 (
    .I(seg_4_2_sp4_v_b_30_15250),
    .O(seg_4_2_local_g3_6_19126)
  );
  LocalMux t2332 (
    .I(seg_4_5_lutff_0_out_15593),
    .O(seg_4_5_local_g1_0_19473)
  );
  LocalMux t2333 (
    .I(seg_5_6_neigh_op_bnl_0_15593),
    .O(seg_5_6_local_g3_0_23443)
  );
  LocalMux t2334 (
    .I(seg_3_5_neigh_op_rgt_3_15596),
    .O(seg_3_5_local_g2_3_15653)
  );
  LocalMux t2335 (
    .I(seg_5_5_neigh_op_lft_3_15596),
    .O(seg_5_5_local_g0_3_23299)
  );
  LocalMux t2336 (
    .I(seg_4_5_lutff_4_out_15597),
    .O(seg_4_5_local_g3_4_19493)
  );
  LocalMux t2337 (
    .I(seg_3_6_neigh_op_bnr_5_15598),
    .O(seg_3_6_local_g1_5_15770)
  );
  LocalMux t2338 (
    .I(seg_4_5_lutff_5_out_15598),
    .O(seg_4_5_local_g1_5_19478)
  );
  LocalMux t2339 (
    .I(seg_4_5_lutff_6_out_15599),
    .O(seg_4_5_local_g1_6_19479)
  );
  CascadeMux t234 (
    .I(net_17169),
    .O(net_17169_cascademuxed)
  );
  LocalMux t2340 (
    .I(seg_5_4_neigh_op_tnl_7_15600),
    .O(seg_5_4_local_g3_7_23204)
  );
  LocalMux t2341 (
    .I(seg_7_5_sp4_h_r_47_19561),
    .O(seg_7_5_local_g2_7_30350)
  );
  LocalMux t2342 (
    .I(seg_7_5_sp4_h_r_9_30432),
    .O(seg_7_5_local_g1_1_30336)
  );
  Span4Mux_h0 t2343 (
    .I(seg_7_5_sp4_h_l_36_15729),
    .O(seg_7_5_sp4_h_r_9_30432)
  );
  LocalMux t2344 (
    .I(seg_9_5_sp4_h_r_27_30426),
    .O(seg_9_5_local_g2_3_38008)
  );
  Span4Mux_h2 t2345 (
    .I(seg_7_5_sp4_h_l_42_15737),
    .O(seg_9_5_sp4_h_r_27_30426)
  );
  LocalMux t2346 (
    .I(seg_7_6_sp4_v_b_44_27237),
    .O(seg_7_6_local_g3_4_30478)
  );
  Span4Mux_v1 t2347 (
    .I(seg_7_5_sp4_h_l_44_15739),
    .O(seg_7_6_sp4_v_b_44_27237)
  );
  LocalMux t2348 (
    .I(seg_5_17_sp4_r_v_b_0_24510),
    .O(seg_5_17_local_g1_0_24780)
  );
  Span4Mux_v4 t2349 (
    .I(seg_6_13_sp4_v_b_4_24022),
    .O(seg_5_17_sp4_r_v_b_0_24510)
  );
  CascadeMux t235 (
    .I(net_17268),
    .O(net_17268_cascademuxed)
  );
  Span4Mux_v4 t2350 (
    .I(seg_6_9_sp4_v_b_4_23530),
    .O(seg_6_13_sp4_v_b_4_24022)
  );
  Span4Mux_v4 t2351 (
    .I(seg_6_5_sp4_h_l_41_11903),
    .O(seg_6_9_sp4_v_b_4_23530)
  );
  LocalMux t2352 (
    .I(seg_16_3_sp4_h_r_11_64655),
    .O(seg_16_3_local_g1_3_64569)
  );
  Span4Mux_h0 t2353 (
    .I(seg_16_3_sp4_h_l_38_49335),
    .O(seg_16_3_sp4_h_r_11_64655)
  );
  Span4Mux_h4 t2354 (
    .I(seg_12_3_sp4_h_l_42_34015),
    .O(seg_16_3_sp4_h_l_38_49335)
  );
  Span4Mux_h4 t2355 (
    .I(seg_8_3_sp4_h_l_41_19319),
    .O(seg_12_3_sp4_h_l_42_34015)
  );
  Span4Mux_h4 t2356 (
    .I(seg_4_3_sp4_v_t_41_15622),
    .O(seg_8_3_sp4_h_l_41_19319)
  );
  LocalMux t2357 (
    .I(seg_4_7_sp4_v_b_18_15746),
    .O(seg_4_7_local_g1_2_19721)
  );
  LocalMux t2358 (
    .I(seg_4_7_sp4_v_b_20_15748),
    .O(seg_4_7_local_g0_4_19715)
  );
  LocalMux t2359 (
    .I(seg_3_6_neigh_op_rgt_0_15716),
    .O(seg_3_6_local_g3_0_15781)
  );
  CascadeMux t236 (
    .I(net_17298),
    .O(net_17298_cascademuxed)
  );
  LocalMux t2360 (
    .I(seg_3_7_neigh_op_bnr_1_15717),
    .O(seg_3_7_local_g1_1_15889)
  );
  LocalMux t2361 (
    .I(seg_3_7_neigh_op_bnr_2_15718),
    .O(seg_3_7_local_g1_2_15890)
  );
  LocalMux t2362 (
    .I(seg_3_7_neigh_op_bnr_3_15719),
    .O(seg_3_7_local_g1_3_15891)
  );
  LocalMux t2363 (
    .I(seg_3_7_neigh_op_bnr_5_15721),
    .O(seg_3_7_local_g0_5_15885)
  );
  LocalMux t2364 (
    .I(seg_3_7_neigh_op_bnr_6_15722),
    .O(seg_3_7_local_g0_6_15886)
  );
  LocalMux t2365 (
    .I(seg_4_6_lutff_7_out_15723),
    .O(seg_4_6_local_g0_7_19595)
  );
  LocalMux t2366 (
    .I(seg_5_16_sp4_v_b_23_20689),
    .O(seg_5_16_local_g0_7_24656)
  );
  Span4Mux_v3 t2367 (
    .I(seg_5_13_sp4_v_b_7_20192),
    .O(seg_5_16_sp4_v_b_23_20689)
  );
  Span4Mux_v4 t2368 (
    .I(seg_5_9_sp4_v_b_4_19699),
    .O(seg_5_13_sp4_v_b_7_20192)
  );
  LocalMux t2369 (
    .I(seg_5_7_neigh_op_lft_1_15840),
    .O(seg_5_7_local_g1_1_23551)
  );
  CascadeMux t237 (
    .I(net_17304),
    .O(net_17304_cascademuxed)
  );
  LocalMux t2370 (
    .I(seg_5_8_neigh_op_bnl_3_15842),
    .O(seg_5_8_local_g2_3_23684)
  );
  LocalMux t2371 (
    .I(seg_5_7_neigh_op_lft_5_15844),
    .O(seg_5_7_local_g1_5_23555)
  );
  LocalMux t2372 (
    .I(seg_4_7_lutff_6_out_15845),
    .O(seg_4_7_local_g1_6_19725)
  );
  LocalMux t2373 (
    .I(seg_4_7_lutff_7_out_15846),
    .O(seg_4_7_local_g0_7_19718)
  );
  LocalMux t2374 (
    .I(seg_4_18_sp4_v_b_14_17095),
    .O(seg_4_18_local_g0_6_21070)
  );
  Span4Mux_v3 t2375 (
    .I(seg_4_15_sp4_v_b_0_16602),
    .O(seg_4_18_sp4_v_b_14_17095)
  );
  Span4Mux_v4 t2376 (
    .I(seg_4_11_sp4_v_b_0_16110),
    .O(seg_4_15_sp4_v_b_0_16602)
  );
  Span4Mux_v4 t2377 (
    .I(seg_4_7_sp4_h_r_0_19805),
    .O(seg_4_11_sp4_v_b_0_16110)
  );
  LocalMux t2378 (
    .I(seg_7_15_sp4_r_v_b_9_31302),
    .O(seg_7_15_local_g2_1_31574)
  );
  Span4Mux_v4 t2379 (
    .I(seg_8_11_sp4_v_b_9_30810),
    .O(seg_7_15_sp4_r_v_b_9_31302)
  );
  CascadeMux t238 (
    .I(net_17421),
    .O(net_17421_cascademuxed)
  );
  Span4Mux_v4 t2380 (
    .I(seg_8_7_sp4_h_l_41_19811),
    .O(seg_8_11_sp4_v_b_9_30810)
  );
  LocalMux t2381 (
    .I(seg_16_3_sp4_h_r_38_53166),
    .O(seg_16_3_local_g2_6_64580)
  );
  Span4Mux_h3 t2382 (
    .I(seg_13_3_sp4_h_l_37_37837),
    .O(seg_16_3_sp4_h_r_38_53166)
  );
  Span4Mux_h4 t2383 (
    .I(seg_9_3_sp4_h_l_44_23155),
    .O(seg_13_3_sp4_h_l_37_37837)
  );
  Span4Mux_h4 t2384 (
    .I(seg_5_3_sp4_v_t_44_19456),
    .O(seg_9_3_sp4_h_l_44_23155)
  );
  LocalMux t2385 (
    .I(seg_2_11_sp4_h_r_23_8345),
    .O(seg_2_11_local_g1_7_12556)
  );
  Span4Mux_h3 t2386 (
    .I(seg_5_11_sp4_v_b_10_19951),
    .O(seg_2_11_sp4_h_r_23_8345)
  );
  LocalMux t2387 (
    .I(seg_2_12_sp4_r_v_b_20_12532),
    .O(seg_2_12_local_g3_4_12692)
  );
  Span4Mux_v3 t2388 (
    .I(seg_3_9_sp4_h_r_3_16225),
    .O(seg_2_12_sp4_r_v_b_20_12532)
  );
  LocalMux t2389 (
    .I(seg_2_11_sp4_r_v_b_27_12526),
    .O(seg_2_11_local_g0_3_12544)
  );
  CascadeMux t239 (
    .I(net_18968),
    .O(net_18968_cascademuxed)
  );
  Span4Mux_v2 t2390 (
    .I(seg_3_9_sp4_h_r_9_16231),
    .O(seg_2_11_sp4_r_v_b_27_12526)
  );
  LocalMux t2391 (
    .I(seg_2_11_sp4_r_v_b_29_12528),
    .O(seg_2_11_local_g1_5_12554)
  );
  Span4Mux_v2 t2392 (
    .I(seg_3_9_sp4_h_r_11_16223),
    .O(seg_2_11_sp4_r_v_b_29_12528)
  );
  LocalMux t2393 (
    .I(seg_2_11_sp4_v_b_24_8209),
    .O(seg_2_11_local_g3_0_12565)
  );
  Span4Mux_v2 t2394 (
    .I(seg_2_9_sp4_h_r_0_12389),
    .O(seg_2_11_sp4_v_b_24_8209)
  );
  LocalMux t2395 (
    .I(seg_2_11_sp4_v_b_26_8211),
    .O(seg_2_11_local_g3_2_12567)
  );
  Span4Mux_v2 t2396 (
    .I(seg_2_9_sp4_h_r_8_12399),
    .O(seg_2_11_sp4_v_b_26_8211)
  );
  LocalMux t2397 (
    .I(seg_2_11_sp4_h_r_21_8353),
    .O(seg_2_11_local_g0_5_12546)
  );
  Span4Mux_h3 t2398 (
    .I(seg_5_11_sp4_v_b_3_19942),
    .O(seg_2_11_sp4_h_r_21_8353)
  );
  LocalMux t2399 (
    .I(seg_2_11_sp4_h_r_16_8350),
    .O(seg_2_11_local_g0_0_12541)
  );
  CascadeMux t24 (
    .I(net_7390),
    .O(net_7390_cascademuxed)
  );
  CascadeMux t240 (
    .I(net_18980),
    .O(net_18980_cascademuxed)
  );
  Span4Mux_h3 t2400 (
    .I(seg_5_11_sp4_v_b_5_19944),
    .O(seg_2_11_sp4_h_r_16_8350)
  );
  LocalMux t2401 (
    .I(seg_2_11_sp4_h_r_17_8349),
    .O(seg_2_11_local_g0_1_12542)
  );
  Span4Mux_h3 t2402 (
    .I(seg_5_11_sp4_v_b_11_19950),
    .O(seg_2_11_sp4_h_r_17_8349)
  );
  LocalMux t2403 (
    .I(seg_2_12_sp4_r_v_b_27_12649),
    .O(seg_2_12_local_g0_3_12667)
  );
  Span4Mux_v2 t2404 (
    .I(seg_3_10_sp4_h_r_9_16354),
    .O(seg_2_12_sp4_r_v_b_27_12649)
  );
  LocalMux t2405 (
    .I(seg_2_12_sp4_r_v_b_29_12651),
    .O(seg_2_12_local_g0_5_12669)
  );
  Span4Mux_v2 t2406 (
    .I(seg_3_10_sp4_h_r_11_16346),
    .O(seg_2_12_sp4_r_v_b_29_12651)
  );
  LocalMux t2407 (
    .I(seg_2_12_sp4_v_b_26_8358),
    .O(seg_2_12_local_g3_2_12690)
  );
  Span4Mux_v2 t2408 (
    .I(seg_2_10_sp4_h_r_2_12516),
    .O(seg_2_12_sp4_v_b_26_8358)
  );
  LocalMux t2409 (
    .I(seg_2_13_sp4_h_r_14_8642),
    .O(seg_2_13_local_g0_6_12793)
  );
  CascadeMux t241 (
    .I(net_18992),
    .O(net_18992_cascademuxed)
  );
  Span4Mux_h3 t2410 (
    .I(seg_5_13_sp4_v_b_10_20197),
    .O(seg_2_13_sp4_h_r_14_8642)
  );
  LocalMux t2411 (
    .I(seg_2_12_sp4_h_r_29_2695),
    .O(seg_2_12_local_g2_5_12685)
  );
  Span4Mux_h2 t2412 (
    .I(seg_4_12_sp4_v_b_0_16233),
    .O(seg_2_12_sp4_h_r_29_2695)
  );
  LocalMux t2413 (
    .I(seg_2_12_sp4_h_r_33_2699),
    .O(seg_2_12_local_g2_1_12681)
  );
  Span4Mux_h2 t2414 (
    .I(seg_4_12_sp4_v_b_4_16237),
    .O(seg_2_12_sp4_h_r_33_2699)
  );
  LocalMux t2415 (
    .I(seg_2_12_sp4_h_r_32_2698),
    .O(seg_2_12_local_g3_0_12688)
  );
  Span4Mux_h2 t2416 (
    .I(seg_4_12_sp4_v_b_8_16241),
    .O(seg_2_12_sp4_h_r_32_2698)
  );
  LocalMux t2417 (
    .I(seg_2_12_sp4_h_r_27_2675),
    .O(seg_2_12_local_g2_3_12683)
  );
  Span4Mux_h2 t2418 (
    .I(seg_4_12_sp4_v_b_10_16243),
    .O(seg_2_12_sp4_h_r_27_2675)
  );
  LocalMux t2419 (
    .I(seg_0_6_sp4_r_v_b_16_1020),
    .O(seg_0_6_local_g3_0_1278)
  );
  CascadeMux t242 (
    .I(net_18998),
    .O(net_18998_cascademuxed)
  );
  Span4Mux_v1 t2420 (
    .I(seg_1_7_sp4_v_t_44_1857),
    .O(seg_0_6_sp4_r_v_b_16_1020)
  );
  Span4Mux_v4 t2421 (
    .I(seg_1_11_sp4_h_r_9_8354),
    .O(seg_1_7_sp4_v_t_44_1857)
  );
  LocalMux t2422 (
    .I(seg_0_24_sp4_r_v_b_19_4884),
    .O(seg_0_24_local_g3_3_5142)
  );
  Span4Mux_v3 t2423 (
    .I(seg_1_21_sp4_h_r_0_9813),
    .O(seg_0_24_sp4_r_v_b_19_4884)
  );
  Span4Mux_h4 t2424 (
    .I(seg_5_21_sp4_v_b_7_21176),
    .O(seg_1_21_sp4_h_r_0_9813)
  );
  Span4Mux_v4 t2425 (
    .I(seg_5_17_sp4_v_b_4_20683),
    .O(seg_5_21_sp4_v_b_7_21176)
  );
  Span4Mux_v4 t2426 (
    .I(seg_5_13_sp4_v_b_1_20186),
    .O(seg_5_17_sp4_v_b_4_20683)
  );
  LocalMux t2427 (
    .I(seg_4_13_sp4_r_v_b_19_20316),
    .O(seg_4_13_local_g3_3_20476)
  );
  LocalMux t2428 (
    .I(seg_0_24_sp4_v_b_10_4446),
    .O(seg_0_24_local_g0_2_5117)
  );
  Span4Mux_v4 t2429 (
    .I(seg_0_20_sp4_v_b_10_3575),
    .O(seg_0_24_sp4_v_b_10_4446)
  );
  CascadeMux t243 (
    .I(net_19004),
    .O(net_19004_cascademuxed)
  );
  Span4Mux_v4 t2430 (
    .I(seg_0_16_sp4_v_b_10_2723),
    .O(seg_0_20_sp4_v_b_10_3575)
  );
  Span4Mux_v4 t2431 (
    .I(seg_0_12_sp4_h_r_4_2686),
    .O(seg_0_16_sp4_v_b_10_2723)
  );
  Span4Mux_h4 t2432 (
    .I(seg_4_12_sp4_v_b_11_16242),
    .O(seg_0_12_sp4_h_r_4_2686)
  );
  LocalMux t2433 (
    .I(seg_0_24_sp4_v_b_19_4669),
    .O(seg_0_24_local_g0_3_5118)
  );
  Span4Mux_v3 t2434 (
    .I(seg_0_21_sp4_h_r_0_4602),
    .O(seg_0_24_sp4_v_b_19_4669)
  );
  Span4Mux_h4 t2435 (
    .I(seg_4_21_sp4_v_b_0_17340),
    .O(seg_0_21_sp4_h_r_0_4602)
  );
  Span4Mux_v4 t2436 (
    .I(seg_4_17_sp4_v_b_0_16848),
    .O(seg_4_21_sp4_v_b_0_17340)
  );
  Span4Mux_v4 t2437 (
    .I(seg_4_13_sp4_v_b_4_16360),
    .O(seg_4_17_sp4_v_b_0_16848)
  );
  LocalMux t2438 (
    .I(seg_4_13_sp4_v_b_6_16362),
    .O(seg_4_13_local_g0_6_20455)
  );
  LocalMux t2439 (
    .I(seg_0_6_sp4_v_b_39_1241),
    .O(seg_0_6_local_g3_7_1285)
  );
  CascadeMux t244 (
    .I(net_19010),
    .O(net_19010_cascademuxed)
  );
  Span4Mux_v3 t2440 (
    .I(seg_0_9_sp4_h_r_2_2040),
    .O(seg_0_6_sp4_v_b_39_1241)
  );
  Span4Mux_h4 t2441 (
    .I(seg_4_9_sp4_v_t_45_16364),
    .O(seg_0_9_sp4_h_r_2_2040)
  );
  LocalMux t2442 (
    .I(seg_0_24_sp4_v_b_21_4671),
    .O(seg_0_24_local_g1_5_5128)
  );
  Span4Mux_v3 t2443 (
    .I(seg_0_21_sp4_v_b_5_3776),
    .O(seg_0_24_sp4_v_b_21_4671)
  );
  Span4Mux_v4 t2444 (
    .I(seg_0_17_sp4_v_b_2_2924),
    .O(seg_0_21_sp4_v_b_5_3776)
  );
  Span4Mux_v4 t2445 (
    .I(seg_0_13_sp4_h_r_8_2907),
    .O(seg_0_17_sp4_v_b_2_2924)
  );
  Span4Mux_h4 t2446 (
    .I(seg_4_13_sp4_v_b_8_16364),
    .O(seg_0_13_sp4_h_r_8_2907)
  );
  LocalMux t2447 (
    .I(seg_4_13_sp4_v_b_10_16366),
    .O(seg_4_13_local_g1_2_20459)
  );
  LocalMux t2448 (
    .I(seg_4_13_sp4_v_b_12_16478),
    .O(seg_4_13_local_g0_4_20453)
  );
  LocalMux t2449 (
    .I(seg_0_6_sp4_v_b_13_802),
    .O(seg_0_6_local_g1_5_1267)
  );
  CascadeMux t245 (
    .I(net_19131),
    .O(net_19131_cascademuxed)
  );
  Span4Mux_v1 t2450 (
    .I(seg_0_7_sp4_h_r_0_1592),
    .O(seg_0_6_sp4_v_b_13_802)
  );
  Span4Mux_h4 t2451 (
    .I(seg_4_7_sp4_v_t_43_16116),
    .O(seg_0_7_sp4_h_r_0_1592)
  );
  LocalMux t2452 (
    .I(seg_0_6_sp4_v_b_12_801),
    .O(seg_0_6_local_g0_4_1258)
  );
  Span4Mux_v1 t2453 (
    .I(seg_0_7_sp4_h_r_8_1638),
    .O(seg_0_6_sp4_v_b_12_801)
  );
  Span4Mux_h4 t2454 (
    .I(seg_4_7_sp4_v_t_45_16118),
    .O(seg_0_7_sp4_h_r_8_1638)
  );
  LocalMux t2455 (
    .I(seg_3_12_neigh_op_rgt_2_16456),
    .O(seg_3_12_local_g2_2_16513)
  );
  LocalMux t2456 (
    .I(seg_7_15_sp4_v_b_18_27949),
    .O(seg_7_15_local_g0_2_31559)
  );
  Span4Mux_v3 t2457 (
    .I(seg_7_12_sp4_h_l_42_16598),
    .O(seg_7_15_sp4_v_b_18_27949)
  );
  LocalMux t2458 (
    .I(seg_3_12_sp4_h_r_13_12758),
    .O(seg_3_12_local_g1_5_16508)
  );
  LocalMux t2459 (
    .I(seg_4_18_sp4_r_v_b_16_20928),
    .O(seg_4_18_local_g3_0_21088)
  );
  CascadeMux t246 (
    .I(net_19137),
    .O(net_19137_cascademuxed)
  );
  Span4Mux_v3 t2460 (
    .I(seg_5_15_sp4_v_b_2_20435),
    .O(seg_4_18_sp4_r_v_b_16_20928)
  );
  LocalMux t2461 (
    .I(seg_3_18_sp4_r_v_b_2_16973),
    .O(seg_3_18_local_g1_2_17243)
  );
  Span4Mux_v4 t2462 (
    .I(seg_4_14_sp4_v_b_2_16481),
    .O(seg_3_18_sp4_r_v_b_2_16973)
  );
  LocalMux t2463 (
    .I(seg_3_18_sp4_r_v_b_4_16975),
    .O(seg_3_18_local_g1_4_17245)
  );
  Span4Mux_v4 t2464 (
    .I(seg_4_14_sp4_v_b_8_16487),
    .O(seg_3_18_sp4_r_v_b_4_16975)
  );
  LocalMux t2465 (
    .I(seg_7_15_sp4_h_r_40_20796),
    .O(seg_7_15_local_g2_0_31573)
  );
  Span4Mux_h3 t2466 (
    .I(seg_4_15_sp4_v_b_11_16611),
    .O(seg_7_15_sp4_h_r_40_20796)
  );
  LocalMux t2467 (
    .I(seg_7_13_sp4_h_r_11_31408),
    .O(seg_7_13_local_g1_3_31322)
  );
  Span4Mux_h0 t2468 (
    .I(seg_7_13_sp4_h_l_38_16717),
    .O(seg_7_13_sp4_h_r_11_31408)
  );
  LocalMux t2469 (
    .I(seg_3_14_neigh_op_rgt_0_16700),
    .O(seg_3_14_local_g2_0_16757)
  );
  CascadeMux t247 (
    .I(net_19143),
    .O(net_19143_cascademuxed)
  );
  LocalMux t2470 (
    .I(seg_3_14_neigh_op_rgt_3_16703),
    .O(seg_3_14_local_g3_3_16768)
  );
  LocalMux t2471 (
    .I(seg_3_15_neigh_op_bnr_3_16703),
    .O(seg_3_15_local_g0_3_16867)
  );
  LocalMux t2472 (
    .I(seg_4_14_lutff_4_out_16704),
    .O(seg_4_14_local_g1_4_20584)
  );
  LocalMux t2473 (
    .I(seg_4_14_lutff_5_out_16705),
    .O(seg_4_14_local_g2_5_20593)
  );
  LocalMux t2474 (
    .I(seg_4_14_lutff_6_out_16706),
    .O(seg_4_14_local_g3_6_20602)
  );
  LocalMux t2475 (
    .I(seg_4_12_sp4_r_v_b_27_20311),
    .O(seg_4_12_local_g1_3_20337)
  );
  LocalMux t2476 (
    .I(seg_4_12_sp4_v_b_38_16603),
    .O(seg_4_12_local_g2_6_20348)
  );
  LocalMux t2477 (
    .I(seg_4_15_lutff_0_out_16823),
    .O(seg_4_15_local_g0_0_20695)
  );
  LocalMux t2478 (
    .I(seg_4_15_lutff_1_out_16824),
    .O(seg_4_15_local_g2_1_20712)
  );
  LocalMux t2479 (
    .I(seg_3_15_neigh_op_rgt_2_16825),
    .O(seg_3_15_local_g3_2_16890)
  );
  CascadeMux t248 (
    .I(net_19149),
    .O(net_19149_cascademuxed)
  );
  LocalMux t2480 (
    .I(seg_3_15_neigh_op_rgt_3_16826),
    .O(seg_3_15_local_g2_3_16883)
  );
  LocalMux t2481 (
    .I(seg_3_15_neigh_op_rgt_4_16827),
    .O(seg_3_15_local_g3_4_16892)
  );
  LocalMux t2482 (
    .I(seg_3_14_neigh_op_tnr_5_16828),
    .O(seg_3_14_local_g3_5_16770)
  );
  LocalMux t2483 (
    .I(seg_4_15_lutff_6_out_16829),
    .O(seg_4_15_local_g3_6_20725)
  );
  LocalMux t2484 (
    .I(seg_4_15_lutff_7_out_16830),
    .O(seg_4_15_local_g3_7_20726)
  );
  LocalMux t2485 (
    .I(seg_4_16_lutff_0_out_16946),
    .O(seg_4_16_local_g0_0_20818)
  );
  LocalMux t2486 (
    .I(seg_3_16_neigh_op_rgt_1_16947),
    .O(seg_3_16_local_g2_1_17004)
  );
  LocalMux t2487 (
    .I(seg_4_16_lutff_4_out_16950),
    .O(seg_4_16_local_g3_4_20846)
  );
  LocalMux t2488 (
    .I(seg_4_16_lutff_5_out_16951),
    .O(seg_4_16_local_g1_5_20831)
  );
  LocalMux t2489 (
    .I(seg_3_15_neigh_op_tnr_6_16952),
    .O(seg_3_15_local_g3_6_16894)
  );
  CascadeMux t249 (
    .I(net_19155),
    .O(net_19155_cascademuxed)
  );
  LocalMux t2490 (
    .I(seg_4_16_lutff_7_out_16953),
    .O(seg_4_16_local_g0_7_20825)
  );
  LocalMux t2491 (
    .I(seg_4_17_lutff_1_out_17070),
    .O(seg_4_17_local_g0_1_20942)
  );
  LocalMux t2492 (
    .I(seg_4_17_lutff_3_out_17072),
    .O(seg_4_17_local_g1_3_20952)
  );
  LocalMux t2493 (
    .I(seg_4_17_lutff_5_out_17074),
    .O(seg_4_17_local_g1_5_20954)
  );
  LocalMux t2494 (
    .I(seg_7_17_sp4_h_r_37_21035),
    .O(seg_7_17_local_g2_5_31824)
  );
  LocalMux t2495 (
    .I(seg_7_17_sp4_h_r_9_31908),
    .O(seg_7_17_local_g1_1_31812)
  );
  Span4Mux_h0 t2496 (
    .I(seg_7_17_sp4_h_l_36_17205),
    .O(seg_7_17_sp4_h_r_9_31908)
  );
  LocalMux t2497 (
    .I(seg_7_17_sp4_h_r_45_21045),
    .O(seg_7_17_local_g3_5_31832)
  );
  LocalMux t2498 (
    .I(seg_5_15_sp4_h_r_7_24629),
    .O(seg_5_15_local_g0_7_24533)
  );
  Span4Mux_h0 t2499 (
    .I(seg_5_15_sp4_v_t_42_20930),
    .O(seg_5_15_sp4_h_r_7_24629)
  );
  CascadeMux t25 (
    .I(net_7402),
    .O(net_7402_cascademuxed)
  );
  CascadeMux t250 (
    .I(net_19161),
    .O(net_19161_cascademuxed)
  );
  LocalMux t2500 (
    .I(seg_4_6_sp4_h_r_10_19684),
    .O(seg_4_6_local_g0_2_19590)
  );
  Span4Mux_h0 t2501 (
    .I(seg_4_6_sp4_v_t_40_15990),
    .O(seg_4_6_sp4_h_r_10_19684)
  );
  Span4Mux_v4 t2502 (
    .I(seg_4_10_sp4_v_t_44_16486),
    .O(seg_4_6_sp4_v_t_40_15990)
  );
  Span4Mux_v4 t2503 (
    .I(seg_4_14_sp4_v_t_43_16977),
    .O(seg_4_10_sp4_v_t_44_16486)
  );
  LocalMux t2504 (
    .I(seg_5_18_neigh_op_tnl_6_17321),
    .O(seg_5_18_local_g3_6_24925)
  );
  LocalMux t2505 (
    .I(seg_4_14_sp4_v_b_27_16726),
    .O(seg_4_14_local_g2_3_20591)
  );
  Span4Mux_v2 t2506 (
    .I(seg_4_16_sp4_v_t_38_17218),
    .O(seg_4_14_sp4_v_b_27_16726)
  );
  LocalMux t2507 (
    .I(seg_4_14_sp4_v_b_32_16733),
    .O(seg_4_14_local_g3_0_20596)
  );
  Span4Mux_v2 t2508 (
    .I(seg_4_16_sp4_v_t_40_17220),
    .O(seg_4_14_sp4_v_b_32_16733)
  );
  LocalMux t2509 (
    .I(seg_5_19_neigh_op_tnl_4_17442),
    .O(seg_5_19_local_g2_4_25038)
  );
  CascadeMux t251 (
    .I(net_19167),
    .O(net_19167_cascademuxed)
  );
  LocalMux t2510 (
    .I(seg_4_19_neigh_op_top_5_17443),
    .O(seg_4_19_local_g0_5_21192)
  );
  LocalMux t2511 (
    .I(seg_4_19_sp4_h_r_1_21282),
    .O(seg_4_19_local_g1_1_21196)
  );
  Span4Mux_h0 t2512 (
    .I(seg_4_19_sp4_v_t_36_17585),
    .O(seg_4_19_sp4_h_r_1_21282)
  );
  LocalMux t2513 (
    .I(seg_3_2_sp4_r_v_b_43_15378),
    .O(seg_3_2_local_g3_3_15292)
  );
  Span4Mux_v3 t2514 (
    .I(seg_4_5_sp4_v_t_47_15874),
    .O(seg_3_2_sp4_r_v_b_43_15378)
  );
  Sp12to4 t2515 (
    .I(seg_4_8_sp12_v_b_23_19804),
    .O(seg_4_5_sp4_v_t_47_15874)
  );
  Span12Mux_v11 t2516 (
    .I(seg_4_19_sp12_v_t_23_21280),
    .O(seg_4_8_sp12_v_b_23_19804)
  );
  LocalMux t2517 (
    .I(seg_4_2_sp4_v_b_47_15382),
    .O(seg_4_2_local_g3_7_19127)
  );
  Span4Mux_v3 t2518 (
    .I(seg_4_5_sp4_v_t_47_15874),
    .O(seg_4_2_sp4_v_b_47_15382)
  );
  LocalMux t2519 (
    .I(seg_4_1_neigh_op_rgt_3_18894),
    .O(seg_4_1_local_g3_3_18960)
  );
  CascadeMux t252 (
    .I(net_19173),
    .O(net_19173_cascademuxed)
  );
  LocalMux t2520 (
    .I(seg_5_1_lutff_3_out_18894),
    .O(seg_5_1_local_g3_3_22791)
  );
  LocalMux t2521 (
    .I(seg_5_0_logic_op_top_7_18898),
    .O(seg_5_0_local_g1_7_22721)
  );
  LocalMux t2522 (
    .I(seg_5_3_neigh_op_bot_5_19024),
    .O(seg_5_3_local_g0_5_23055)
  );
  LocalMux t2523 (
    .I(seg_8_3_sp4_h_r_30_26919),
    .O(seg_8_3_local_g2_6_33934)
  );
  Span4Mux_h2 t2524 (
    .I(seg_6_3_sp4_v_b_6_22898),
    .O(seg_8_3_sp4_h_r_30_26919)
  );
  LocalMux t2525 (
    .I(seg_6_3_neigh_op_lft_2_19180),
    .O(seg_6_3_local_g0_2_26839)
  );
  LocalMux t2526 (
    .I(seg_6_3_neigh_op_lft_2_19180),
    .O(seg_6_3_local_g1_2_26847)
  );
  LocalMux t2527 (
    .I(seg_6_4_neigh_op_bnl_2_19180),
    .O(seg_6_4_local_g2_2_26957)
  );
  LocalMux t2528 (
    .I(seg_6_4_neigh_op_bnl_2_19180),
    .O(seg_6_4_local_g3_2_26965)
  );
  LocalMux t2529 (
    .I(seg_5_3_lutff_5_out_19183),
    .O(seg_5_3_local_g2_5_23071)
  );
  CascadeMux t253 (
    .I(net_19254),
    .O(net_19254_cascademuxed)
  );
  LocalMux t2530 (
    .I(seg_5_16_sp4_v_b_13_20679),
    .O(seg_5_16_local_g0_5_24654)
  );
  Span4Mux_v3 t2531 (
    .I(seg_5_13_sp4_v_b_9_20194),
    .O(seg_5_16_sp4_v_b_13_20679)
  );
  Span4Mux_v4 t2532 (
    .I(seg_5_9_sp4_v_b_9_19702),
    .O(seg_5_13_sp4_v_b_9_20194)
  );
  Span4Mux_v4 t2533 (
    .I(seg_5_5_sp4_v_b_6_19209),
    .O(seg_5_9_sp4_v_b_9_19702)
  );
  LocalMux t2534 (
    .I(seg_5_7_sp4_v_b_4_19453),
    .O(seg_5_7_local_g1_4_23554)
  );
  Span4Mux_v4 t2535 (
    .I(seg_5_3_sp4_v_b_8_19069),
    .O(seg_5_7_sp4_v_b_4_19453)
  );
  LocalMux t2536 (
    .I(seg_4_5_neigh_op_bnr_6_19307),
    .O(seg_4_5_local_g0_6_19471)
  );
  LocalMux t2537 (
    .I(seg_8_4_sp4_h_r_11_34132),
    .O(seg_8_4_local_g0_3_34038)
  );
  Span4Mux_h0 t2538 (
    .I(seg_8_4_sp4_h_l_38_19441),
    .O(seg_8_4_sp4_h_r_11_34132)
  );
  LocalMux t2539 (
    .I(seg_7_4_sp4_h_r_28_23273),
    .O(seg_7_4_local_g3_4_30232)
  );
  CascadeMux t254 (
    .I(net_19260),
    .O(net_19260_cascademuxed)
  );
  LocalMux t2540 (
    .I(seg_5_6_sp4_r_v_b_19_23286),
    .O(seg_5_6_local_g3_3_23446)
  );
  LocalMux t2541 (
    .I(seg_5_6_sp4_r_v_b_21_23288),
    .O(seg_5_6_local_g3_5_23448)
  );
  LocalMux t2542 (
    .I(seg_5_6_sp4_v_b_0_19326),
    .O(seg_5_6_local_g0_0_23419)
  );
  LocalMux t2543 (
    .I(seg_5_6_sp4_v_b_8_19334),
    .O(seg_5_6_local_g1_0_23427)
  );
  LocalMux t2544 (
    .I(seg_5_6_sp4_v_b_10_19336),
    .O(seg_5_6_local_g0_2_23421)
  );
  LocalMux t2545 (
    .I(seg_5_6_sp4_v_b_12_19448),
    .O(seg_5_6_local_g0_4_23423)
  );
  LocalMux t2546 (
    .I(seg_5_6_sp4_v_b_14_19450),
    .O(seg_5_6_local_g0_6_23425)
  );
  LocalMux t2547 (
    .I(seg_4_5_neigh_op_rgt_7_19431),
    .O(seg_4_5_local_g2_7_19488)
  );
  LocalMux t2548 (
    .I(seg_8_5_sp4_h_r_47_23392),
    .O(seg_8_5_local_g2_7_34181)
  );
  LocalMux t2549 (
    .I(seg_3_5_sp4_h_r_10_15730),
    .O(seg_3_5_local_g1_2_15644)
  );
  CascadeMux t255 (
    .I(net_19266),
    .O(net_19266_cascademuxed)
  );
  LocalMux t2550 (
    .I(seg_3_5_sp4_h_r_12_11898),
    .O(seg_3_5_local_g0_4_15638)
  );
  LocalMux t2551 (
    .I(seg_3_5_sp4_h_r_14_11902),
    .O(seg_3_5_local_g0_6_15640)
  );
  LocalMux t2552 (
    .I(seg_2_5_sp4_h_r_5_11904),
    .O(seg_2_5_local_g1_5_11816)
  );
  LocalMux t2553 (
    .I(seg_7_6_sp4_h_r_13_27217),
    .O(seg_7_6_local_g0_5_30455)
  );
  Span4Mux_h1 t2554 (
    .I(seg_6_6_sp4_v_b_0_23157),
    .O(seg_7_6_sp4_h_r_13_27217)
  );
  LocalMux t2555 (
    .I(seg_5_5_neigh_op_top_1_19548),
    .O(seg_5_5_local_g1_1_23305)
  );
  LocalMux t2556 (
    .I(seg_5_5_neigh_op_top_2_19549),
    .O(seg_5_5_local_g1_2_23306)
  );
  LocalMux t2557 (
    .I(seg_5_5_neigh_op_top_3_19550),
    .O(seg_5_5_local_g1_3_23307)
  );
  LocalMux t2558 (
    .I(seg_5_5_neigh_op_top_4_19551),
    .O(seg_5_5_local_g1_4_23308)
  );
  LocalMux t2559 (
    .I(seg_5_5_neigh_op_top_5_19552),
    .O(seg_5_5_local_g0_5_23301)
  );
  CascadeMux t256 (
    .I(net_19272),
    .O(net_19272_cascademuxed)
  );
  LocalMux t2560 (
    .I(seg_5_5_neigh_op_top_6_19553),
    .O(seg_5_5_local_g1_6_23310)
  );
  LocalMux t2561 (
    .I(seg_15_6_sp4_h_r_8_61200),
    .O(seg_15_6_local_g1_0_61104)
  );
  Span4Mux_h0 t2562 (
    .I(seg_15_6_sp4_h_l_40_45875),
    .O(seg_15_6_sp4_h_r_8_61200)
  );
  Span4Mux_h4 t2563 (
    .I(seg_11_6_sp4_h_l_39_30548),
    .O(seg_15_6_sp4_h_l_40_45875)
  );
  Span4Mux_h4 t2564 (
    .I(seg_7_6_sp4_h_l_43_15859),
    .O(seg_11_6_sp4_h_l_39_30548)
  );
  LocalMux t2565 (
    .I(seg_4_7_neigh_op_rgt_3_19673),
    .O(seg_4_7_local_g3_3_19738)
  );
  LocalMux t2566 (
    .I(seg_5_8_neigh_op_bot_3_19673),
    .O(seg_5_8_local_g1_3_23676)
  );
  LocalMux t2567 (
    .I(seg_5_16_sp12_v_b_3_23389),
    .O(seg_5_16_local_g3_3_24676)
  );
  LocalMux t2568 (
    .I(seg_7_15_sp4_r_v_b_3_31296),
    .O(seg_7_15_local_g1_3_31568)
  );
  Span4Mux_v4 t2569 (
    .I(seg_8_11_sp4_v_b_0_30803),
    .O(seg_7_15_sp4_r_v_b_3_31296)
  );
  CascadeMux t257 (
    .I(net_19284),
    .O(net_19284_cascademuxed)
  );
  Span4Mux_v4 t2570 (
    .I(seg_8_7_sp4_h_l_42_19814),
    .O(seg_8_11_sp4_v_b_0_30803)
  );
  LocalMux t2571 (
    .I(seg_7_15_sp4_h_r_23_28137),
    .O(seg_7_15_local_g1_7_31572)
  );
  Span4Mux_h1 t2572 (
    .I(seg_6_15_sp4_v_b_10_24274),
    .O(seg_7_15_sp4_h_r_23_28137)
  );
  Span4Mux_v4 t2573 (
    .I(seg_6_11_sp4_v_b_7_23777),
    .O(seg_6_15_sp4_v_b_10_24274)
  );
  Span4Mux_v4 t2574 (
    .I(seg_6_7_sp4_v_b_11_23289),
    .O(seg_6_11_sp4_v_b_7_23777)
  );
  LocalMux t2575 (
    .I(seg_5_7_neigh_op_top_3_19796),
    .O(seg_5_7_local_g1_3_23553)
  );
  LocalMux t2576 (
    .I(seg_5_8_lutff_5_out_19798),
    .O(seg_5_8_local_g1_5_23678)
  );
  LocalMux t2577 (
    .I(seg_5_8_lutff_6_out_19799),
    .O(seg_5_8_local_g2_6_23687)
  );
  LocalMux t2578 (
    .I(seg_7_8_sp4_h_r_38_19933),
    .O(seg_7_8_local_g2_6_30718)
  );
  LocalMux t2579 (
    .I(seg_7_8_sp4_h_r_44_19939),
    .O(seg_7_8_local_g3_4_30724)
  );
  CascadeMux t258 (
    .I(net_19290),
    .O(net_19290_cascademuxed)
  );
  LocalMux t2580 (
    .I(seg_9_11_sp4_v_b_19_34763),
    .O(seg_9_11_local_g1_3_38738)
  );
  Span4Mux_v3 t2581 (
    .I(seg_9_8_sp4_h_l_43_23767),
    .O(seg_9_11_sp4_v_b_19_34763)
  );
  LocalMux t2582 (
    .I(seg_7_8_sp4_h_r_32_23769),
    .O(seg_7_8_local_g2_0_30712)
  );
  LocalMux t2583 (
    .I(seg_7_4_sp4_h_r_12_27014),
    .O(seg_7_4_local_g0_4_30208)
  );
  Span4Mux_h1 t2584 (
    .I(seg_6_4_sp4_v_t_36_23402),
    .O(seg_7_4_sp4_h_r_12_27014)
  );
  LocalMux t2585 (
    .I(seg_4_5_sp4_h_r_34_11899),
    .O(seg_4_5_local_g2_2_19483)
  );
  Span4Mux_h2 t2586 (
    .I(seg_6_5_sp4_v_t_47_23536),
    .O(seg_4_5_sp4_h_r_34_11899)
  );
  LocalMux t2587 (
    .I(seg_7_5_sp4_h_r_14_27120),
    .O(seg_7_5_local_g1_6_30341)
  );
  Span4Mux_h1 t2588 (
    .I(seg_6_5_sp4_v_t_47_23536),
    .O(seg_7_5_sp4_h_r_14_27120)
  );
  LocalMux t2589 (
    .I(seg_5_6_sp4_v_b_26_19574),
    .O(seg_5_6_local_g3_2_23445)
  );
  CascadeMux t259 (
    .I(net_19296),
    .O(net_19296_cascademuxed)
  );
  LocalMux t2590 (
    .I(seg_0_16_sp12_v_b_10_2014),
    .O(seg_0_16_local_g2_2_3392)
  );
  Span12Mux_v7 t2591 (
    .I(seg_0_9_sp12_h_r_1_1991),
    .O(seg_0_16_sp12_v_b_10_2014)
  );
  LocalMux t2592 (
    .I(seg_0_16_sp4_v_b_23_2932),
    .O(seg_0_16_local_g1_7_3389)
  );
  Span4Mux_v3 t2593 (
    .I(seg_0_13_sp4_h_r_4_2895),
    .O(seg_0_16_sp4_v_b_23_2932)
  );
  Span4Mux_h4 t2594 (
    .I(seg_4_13_sp4_v_b_11_16365),
    .O(seg_0_13_sp4_h_r_4_2895)
  );
  Span4Mux_v4 t2595 (
    .I(seg_4_9_sp4_h_r_5_20058),
    .O(seg_4_13_sp4_v_b_11_16365)
  );
  LocalMux t2596 (
    .I(seg_0_11_sp4_v_b_33_2096),
    .O(seg_0_11_local_g2_1_2331)
  );
  Span4Mux_v2 t2597 (
    .I(seg_0_9_sp4_h_r_9_2075),
    .O(seg_0_11_sp4_v_b_33_2096)
  );
  Span4Mux_h4 t2598 (
    .I(seg_4_9_sp4_h_r_9_20062),
    .O(seg_0_9_sp4_h_r_9_2075)
  );
  LocalMux t2599 (
    .I(seg_0_11_sp4_v_b_29_2092),
    .O(seg_0_11_local_g3_5_2343)
  );
  CascadeMux t26 (
    .I(net_7408),
    .O(net_7408_cascademuxed)
  );
  CascadeMux t260 (
    .I(net_19377),
    .O(net_19377_cascademuxed)
  );
  Span4Mux_v2 t2600 (
    .I(seg_0_9_sp4_h_r_11_2031),
    .O(seg_0_11_sp4_v_b_29_2092)
  );
  Span4Mux_h4 t2601 (
    .I(seg_4_9_sp4_h_r_11_20054),
    .O(seg_0_9_sp4_h_r_11_2031)
  );
  LocalMux t2602 (
    .I(seg_0_11_sp4_h_r_26_2463),
    .O(seg_0_11_local_g3_2_2340)
  );
  Span4Mux_h2 t2603 (
    .I(seg_2_11_sp4_h_r_6_12643),
    .O(seg_0_11_sp4_h_r_26_2463)
  );
  Span4Mux_h4 t2604 (
    .I(seg_6_11_sp4_v_b_1_23771),
    .O(seg_2_11_sp4_h_r_6_12643)
  );
  LocalMux t2605 (
    .I(seg_0_11_sp4_h_r_35_2473),
    .O(seg_0_11_local_g2_3_2333)
  );
  Span4Mux_h2 t2606 (
    .I(seg_2_11_sp4_h_r_8_12645),
    .O(seg_0_11_sp4_h_r_35_2473)
  );
  Span4Mux_h4 t2607 (
    .I(seg_6_11_sp4_v_b_3_23773),
    .O(seg_2_11_sp4_h_r_8_12645)
  );
  LocalMux t2608 (
    .I(seg_0_11_sp4_h_r_30_2468),
    .O(seg_0_11_local_g2_6_2336)
  );
  Span4Mux_h2 t2609 (
    .I(seg_2_11_sp4_h_r_10_12637),
    .O(seg_0_11_sp4_h_r_30_2468)
  );
  CascadeMux t261 (
    .I(net_19395),
    .O(net_19395_cascademuxed)
  );
  Span4Mux_h4 t2610 (
    .I(seg_6_11_sp4_v_b_5_23775),
    .O(seg_2_11_sp4_h_r_10_12637)
  );
  LocalMux t2611 (
    .I(seg_0_11_sp4_h_r_33_2471),
    .O(seg_0_11_local_g3_1_2339)
  );
  Span4Mux_h2 t2612 (
    .I(seg_2_11_sp4_h_r_9_12646),
    .O(seg_0_11_sp4_h_r_33_2471)
  );
  Span4Mux_h4 t2613 (
    .I(seg_6_11_sp4_v_b_9_23779),
    .O(seg_2_11_sp4_h_r_9_12646)
  );
  LocalMux t2614 (
    .I(seg_0_11_sp4_h_r_31_2469),
    .O(seg_0_11_local_g3_7_2345)
  );
  Span4Mux_h2 t2615 (
    .I(seg_2_11_sp4_h_r_4_12641),
    .O(seg_0_11_sp4_h_r_31_2469)
  );
  Span4Mux_h4 t2616 (
    .I(seg_6_11_sp4_v_b_11_23781),
    .O(seg_2_11_sp4_h_r_4_12641)
  );
  LocalMux t2617 (
    .I(seg_0_16_sp4_r_v_b_0_2910),
    .O(seg_0_16_local_g1_0_3382)
  );
  Span4Mux_v4 t2618 (
    .I(seg_1_12_sp4_h_r_6_8498),
    .O(seg_0_16_sp4_r_v_b_0_2910)
  );
  Span4Mux_h4 t2619 (
    .I(seg_5_12_sp4_v_b_1_20063),
    .O(seg_1_12_sp4_h_r_6_8498)
  );
  CascadeMux t262 (
    .I(net_19401),
    .O(net_19401_cascademuxed)
  );
  LocalMux t2620 (
    .I(seg_0_16_sp4_r_v_b_8_2918),
    .O(seg_0_16_local_g2_0_3390)
  );
  Span4Mux_v4 t2621 (
    .I(seg_1_12_sp4_h_r_8_8500),
    .O(seg_0_16_sp4_r_v_b_8_2918)
  );
  Span4Mux_h4 t2622 (
    .I(seg_5_12_sp4_v_b_3_20065),
    .O(seg_1_12_sp4_h_r_8_8500)
  );
  LocalMux t2623 (
    .I(seg_0_16_sp4_r_v_b_11_2919),
    .O(seg_0_16_local_g2_3_3393)
  );
  Span4Mux_v4 t2624 (
    .I(seg_1_12_sp4_h_r_5_8497),
    .O(seg_0_16_sp4_r_v_b_11_2919)
  );
  Span4Mux_h4 t2625 (
    .I(seg_5_12_sp4_v_b_5_20067),
    .O(seg_1_12_sp4_h_r_5_8497)
  );
  LocalMux t2626 (
    .I(seg_0_16_sp4_h_r_45_3544),
    .O(seg_0_16_local_g2_5_3395)
  );
  Span4Mux_h1 t2627 (
    .I(seg_1_16_sp4_h_r_8_9088),
    .O(seg_0_16_sp4_h_r_45_3544)
  );
  Span4Mux_h4 t2628 (
    .I(seg_5_16_sp4_v_b_3_20557),
    .O(seg_1_16_sp4_h_r_8_9088)
  );
  Span4Mux_v4 t2629 (
    .I(seg_5_12_sp4_v_b_7_20069),
    .O(seg_5_16_sp4_v_b_3_20557)
  );
  CascadeMux t263 (
    .I(net_19413),
    .O(net_19413_cascademuxed)
  );
  LocalMux t2630 (
    .I(seg_0_16_sp4_r_v_b_3_2911),
    .O(seg_0_16_local_g1_3_3385)
  );
  Span4Mux_v4 t2631 (
    .I(seg_1_12_sp4_h_r_9_8501),
    .O(seg_0_16_sp4_r_v_b_3_2911)
  );
  Span4Mux_h4 t2632 (
    .I(seg_5_12_sp4_v_b_9_20071),
    .O(seg_1_12_sp4_h_r_9_8501)
  );
  LocalMux t2633 (
    .I(seg_0_11_sp4_r_v_b_16_2080),
    .O(seg_0_11_local_g3_0_2338)
  );
  Span4Mux_v3 t2634 (
    .I(seg_1_8_sp4_h_r_5_7909),
    .O(seg_0_11_sp4_r_v_b_16_2080)
  );
  Span4Mux_h4 t2635 (
    .I(seg_5_8_sp4_v_t_46_20073),
    .O(seg_1_8_sp4_h_r_5_7909)
  );
  LocalMux t2636 (
    .I(seg_0_16_sp4_r_v_b_4_2914),
    .O(seg_0_16_local_g1_4_3386)
  );
  Span4Mux_v4 t2637 (
    .I(seg_1_12_sp4_h_r_4_8496),
    .O(seg_0_16_sp4_r_v_b_4_2914)
  );
  Span4Mux_h4 t2638 (
    .I(seg_5_12_sp4_v_b_11_20073),
    .O(seg_1_12_sp4_h_r_4_8496)
  );
  LocalMux t2639 (
    .I(seg_5_16_sp12_v_b_0_23266),
    .O(seg_5_16_local_g2_0_24665)
  );
  LocalMux t2640 (
    .I(seg_4_18_sp4_r_v_b_6_20808),
    .O(seg_4_18_local_g1_6_21078)
  );
  Span4Mux_v4 t2641 (
    .I(seg_5_14_sp4_v_b_10_20320),
    .O(seg_4_18_sp4_r_v_b_6_20808)
  );
  Span4Mux_v4 t2642 (
    .I(seg_5_10_sp4_h_r_10_24007),
    .O(seg_5_14_sp4_v_b_10_20320)
  );
  LocalMux t2643 (
    .I(seg_3_18_sp4_r_v_b_8_16979),
    .O(seg_3_18_local_g2_0_17249)
  );
  Span4Mux_v4 t2644 (
    .I(seg_4_14_sp4_v_b_5_16482),
    .O(seg_3_18_sp4_r_v_b_8_16979)
  );
  Span4Mux_v4 t2645 (
    .I(seg_4_10_sp4_h_r_5_20181),
    .O(seg_4_14_sp4_v_b_5_16482)
  );
  LocalMux t2646 (
    .I(seg_7_15_sp4_h_r_16_28142),
    .O(seg_7_15_local_g1_0_31565)
  );
  Span4Mux_h1 t2647 (
    .I(seg_6_15_sp4_v_b_5_24267),
    .O(seg_7_15_sp4_h_r_16_28142)
  );
  Span4Mux_v4 t2648 (
    .I(seg_6_11_sp4_v_b_2_23774),
    .O(seg_6_15_sp4_v_b_5_24267)
  );
  LocalMux t2649 (
    .I(seg_7_15_sp4_h_r_21_28145),
    .O(seg_7_15_local_g0_5_31562)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t265 (
    .carryinitin(),
    .carryinitout(t264)
  );
  Span4Mux_h1 t2650 (
    .I(seg_6_15_sp4_v_b_2_24266),
    .O(seg_7_15_sp4_h_r_21_28145)
  );
  Span4Mux_v4 t2651 (
    .I(seg_6_11_sp4_v_b_6_23778),
    .O(seg_6_15_sp4_v_b_2_24266)
  );
  LocalMux t2652 (
    .I(seg_5_16_sp4_r_v_b_23_24520),
    .O(seg_5_16_local_g3_7_24680)
  );
  Span4Mux_v3 t2653 (
    .I(seg_6_13_sp4_v_b_2_24020),
    .O(seg_5_16_sp4_r_v_b_23_24520)
  );
  LocalMux t2654 (
    .I(seg_7_15_sp4_h_r_29_24627),
    .O(seg_7_15_local_g2_5_31578)
  );
  Span4Mux_h2 t2655 (
    .I(seg_5_15_sp4_v_b_5_20436),
    .O(seg_7_15_sp4_h_r_29_24627)
  );
  Span4Mux_v4 t2656 (
    .I(seg_5_11_sp4_v_b_9_19948),
    .O(seg_5_15_sp4_v_b_5_20436)
  );
  LocalMux t2657 (
    .I(seg_5_16_sp4_v_b_16_20682),
    .O(seg_5_16_local_g0_0_24649)
  );
  Span4Mux_v3 t2658 (
    .I(seg_5_13_sp4_v_b_5_20190),
    .O(seg_5_16_sp4_v_b_16_20682)
  );
  LocalMux t2659 (
    .I(seg_7_11_sp4_h_r_42_20306),
    .O(seg_7_11_local_g3_2_31091)
  );
  CascadeMux t266 (
    .I(net_19500),
    .O(net_19500_cascademuxed)
  );
  LocalMux t2660 (
    .I(seg_0_11_sp4_h_r_17_2453),
    .O(seg_0_11_local_g0_1_2315)
  );
  Span4Mux_h3 t2661 (
    .I(seg_3_11_sp4_h_r_8_16476),
    .O(seg_0_11_sp4_h_r_17_2453)
  );
  LocalMux t2662 (
    .I(seg_7_11_sp4_h_r_30_24136),
    .O(seg_7_11_local_g3_6_31095)
  );
  LocalMux t2663 (
    .I(seg_0_6_sp4_r_v_b_43_1439),
    .O(seg_0_6_local_g3_3_1281)
  );
  Span4Mux_v3 t2664 (
    .I(seg_1_9_sp4_h_r_6_8057),
    .O(seg_0_6_sp4_r_v_b_43_1439)
  );
  Span4Mux_h4 t2665 (
    .I(seg_5_9_sp4_v_t_37_20187),
    .O(seg_1_9_sp4_h_r_6_8057)
  );
  LocalMux t2666 (
    .I(seg_0_24_sp4_r_v_b_17_4882),
    .O(seg_0_24_local_g3_1_5140)
  );
  Span4Mux_v3 t2667 (
    .I(seg_1_21_sp4_v_b_8_3978),
    .O(seg_0_24_sp4_r_v_b_17_4882)
  );
  Span4Mux_v4 t2668 (
    .I(seg_1_17_sp4_v_b_5_3140),
    .O(seg_1_21_sp4_v_b_8_3978)
  );
  Span4Mux_v4 t2669 (
    .I(seg_1_13_sp4_h_r_5_8644),
    .O(seg_1_17_sp4_v_b_5_3140)
  );
  CascadeMux t267 (
    .I(net_19524),
    .O(net_19524_cascademuxed)
  );
  Span4Mux_h4 t2670 (
    .I(seg_5_13_sp4_v_b_0_20187),
    .O(seg_1_13_sp4_h_r_5_8644)
  );
  LocalMux t2671 (
    .I(seg_0_6_sp4_r_v_b_36_1432),
    .O(seg_0_6_local_g2_4_1274)
  );
  Span4Mux_v3 t2672 (
    .I(seg_1_9_sp4_h_r_8_8059),
    .O(seg_0_6_sp4_r_v_b_36_1432)
  );
  Span4Mux_h4 t2673 (
    .I(seg_5_9_sp4_v_t_39_20189),
    .O(seg_1_9_sp4_h_r_8_8059)
  );
  LocalMux t2674 (
    .I(seg_0_24_sp4_r_v_b_23_4888),
    .O(seg_0_24_local_g3_7_5146)
  );
  Span4Mux_v3 t2675 (
    .I(seg_1_21_sp4_h_r_10_9815),
    .O(seg_0_24_sp4_r_v_b_23_4888)
  );
  Span4Mux_h4 t2676 (
    .I(seg_5_21_sp4_v_b_5_21174),
    .O(seg_1_21_sp4_h_r_10_9815)
  );
  Span4Mux_v4 t2677 (
    .I(seg_5_17_sp4_v_b_2_20681),
    .O(seg_5_21_sp4_v_b_5_21174)
  );
  Span4Mux_v4 t2678 (
    .I(seg_5_13_sp4_v_b_2_20189),
    .O(seg_5_17_sp4_v_b_2_20681)
  );
  LocalMux t2679 (
    .I(seg_0_6_sp4_r_v_b_41_1437),
    .O(seg_0_6_local_g3_1_1279)
  );
  CascadeMux t268 (
    .I(net_19530),
    .O(net_19530_cascademuxed)
  );
  Span4Mux_v3 t2680 (
    .I(seg_1_9_sp4_h_r_4_8055),
    .O(seg_0_6_sp4_r_v_b_41_1437)
  );
  Span4Mux_h4 t2681 (
    .I(seg_5_9_sp4_v_t_41_20191),
    .O(seg_1_9_sp4_h_r_4_8055)
  );
  LocalMux t2682 (
    .I(seg_0_24_sp4_r_v_b_21_4886),
    .O(seg_0_24_local_g3_5_5144)
  );
  Span4Mux_v3 t2683 (
    .I(seg_1_21_sp4_h_r_8_9823),
    .O(seg_0_24_sp4_r_v_b_21_4886)
  );
  Span4Mux_h4 t2684 (
    .I(seg_5_21_sp4_v_b_3_21172),
    .O(seg_1_21_sp4_h_r_8_9823)
  );
  Span4Mux_v4 t2685 (
    .I(seg_5_17_sp4_v_b_7_20684),
    .O(seg_5_21_sp4_v_b_3_21172)
  );
  Span4Mux_v4 t2686 (
    .I(seg_5_13_sp4_v_b_4_20191),
    .O(seg_5_17_sp4_v_b_7_20684)
  );
  LocalMux t2687 (
    .I(seg_0_16_sp4_r_v_b_18_3142),
    .O(seg_0_16_local_g3_2_3400)
  );
  Span4Mux_v3 t2688 (
    .I(seg_1_13_sp4_h_r_1_8638),
    .O(seg_0_16_sp4_r_v_b_18_3142)
  );
  Span4Mux_h4 t2689 (
    .I(seg_5_13_sp4_v_b_8_20195),
    .O(seg_1_13_sp4_h_r_1_8638)
  );
  CascadeMux t269 (
    .I(net_19536),
    .O(net_19536_cascademuxed)
  );
  LocalMux t2690 (
    .I(seg_0_24_sp4_r_v_b_27_5089),
    .O(seg_0_24_local_g1_3_5126)
  );
  Span4Mux_v2 t2691 (
    .I(seg_1_22_sp4_v_b_7_4202),
    .O(seg_0_24_sp4_r_v_b_27_5089)
  );
  Span4Mux_v4 t2692 (
    .I(seg_1_18_sp4_h_r_1_9373),
    .O(seg_1_22_sp4_v_b_7_4202)
  );
  Span4Mux_h4 t2693 (
    .I(seg_5_18_sp4_v_b_1_20801),
    .O(seg_1_18_sp4_h_r_1_9373)
  );
  Span4Mux_v4 t2694 (
    .I(seg_5_14_sp4_v_b_1_20309),
    .O(seg_5_18_sp4_v_b_1_20801)
  );
  LocalMux t2695 (
    .I(seg_0_6_sp4_r_v_b_14_1018),
    .O(seg_0_6_local_g2_6_1276)
  );
  Span4Mux_v1 t2696 (
    .I(seg_1_7_sp4_h_r_10_7757),
    .O(seg_0_6_sp4_r_v_b_14_1018)
  );
  Span4Mux_h4 t2697 (
    .I(seg_5_7_sp4_v_t_41_19945),
    .O(seg_1_7_sp4_h_r_10_7757)
  );
  LocalMux t2698 (
    .I(seg_0_6_sp4_h_r_42_1421),
    .O(seg_0_6_local_g2_2_1272)
  );
  Span4Mux_h1 t2699 (
    .I(seg_1_6_sp4_h_r_7_7617),
    .O(seg_0_6_sp4_h_r_42_1421)
  );
  CascadeMux t27 (
    .I(net_7543),
    .O(net_7543_cascademuxed)
  );
  Span4Mux_h4 t2700 (
    .I(seg_5_6_sp4_v_t_42_19823),
    .O(seg_1_6_sp4_h_r_7_7617)
  );
  Span4Mux_v4 t2701 (
    .I(seg_5_10_sp4_v_t_46_20319),
    .O(seg_5_6_sp4_v_t_42_19823)
  );
  LocalMux t2702 (
    .I(seg_0_24_sp4_r_v_b_34_5098),
    .O(seg_0_24_local_g2_2_5133)
  );
  Span4Mux_v2 t2703 (
    .I(seg_1_22_sp4_v_b_2_4199),
    .O(seg_0_24_sp4_r_v_b_34_5098)
  );
  Span4Mux_v4 t2704 (
    .I(seg_1_18_sp4_h_r_2_9376),
    .O(seg_1_22_sp4_v_b_2_4199)
  );
  Span4Mux_h4 t2705 (
    .I(seg_5_18_sp4_v_b_2_20804),
    .O(seg_1_18_sp4_h_r_2_9376)
  );
  Span4Mux_v4 t2706 (
    .I(seg_5_14_sp4_v_b_11_20319),
    .O(seg_5_18_sp4_v_b_2_20804)
  );
  LocalMux t2707 (
    .I(seg_5_12_lutff_2_out_20287),
    .O(seg_5_12_local_g2_2_24175)
  );
  LocalMux t2708 (
    .I(seg_5_12_lutff_4_out_20289),
    .O(seg_5_12_local_g2_4_24177)
  );
  LocalMux t2709 (
    .I(seg_5_2_sp12_v_b_20_22746),
    .O(seg_5_2_local_g3_4_22955)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t271 (
    .carryinitin(),
    .carryinitout(t270)
  );
  LocalMux t2710 (
    .I(seg_5_3_sp12_v_b_19_22746),
    .O(seg_5_3_local_g2_3_23069)
  );
  LocalMux t2711 (
    .I(seg_5_10_sp12_v_b_4_22746),
    .O(seg_5_10_local_g3_4_23939)
  );
  LocalMux t2712 (
    .I(seg_16_10_sp4_v_b_33_61579),
    .O(seg_16_10_local_g3_1_65444)
  );
  Span4Mux_v2 t2713 (
    .I(seg_16_12_sp4_h_l_38_50442),
    .O(seg_16_10_sp4_v_b_33_61579)
  );
  Span4Mux_h4 t2714 (
    .I(seg_12_12_sp4_h_l_38_35118),
    .O(seg_16_12_sp4_h_l_38_50442)
  );
  Span4Mux_h4 t2715 (
    .I(seg_8_12_sp4_h_l_42_20429),
    .O(seg_12_12_sp4_h_l_38_35118)
  );
  LocalMux t2716 (
    .I(seg_8_6_sp4_v_b_31_30439),
    .O(seg_8_6_local_g2_7_34304)
  );
  Span4Mux_v2 t2717 (
    .I(seg_8_8_sp4_v_t_46_30935),
    .O(seg_8_6_sp4_v_b_31_30439)
  );
  Span4Mux_v4 t2718 (
    .I(seg_8_12_sp4_h_l_46_20423),
    .O(seg_8_8_sp4_v_t_46_30935)
  );
  LocalMux t2719 (
    .I(seg_8_7_sp4_v_b_18_30439),
    .O(seg_8_7_local_g0_2_34406)
  );
  CascadeMux t272 (
    .I(net_19623),
    .O(net_19623_cascademuxed)
  );
  Span4Mux_v1 t2720 (
    .I(seg_8_8_sp4_v_t_46_30935),
    .O(seg_8_7_sp4_v_b_18_30439)
  );
  LocalMux t2721 (
    .I(seg_16_10_sp4_v_b_35_61581),
    .O(seg_16_10_local_g2_3_65438)
  );
  Span4Mux_v2 t2722 (
    .I(seg_16_12_sp4_h_l_46_50440),
    .O(seg_16_10_sp4_v_b_35_61581)
  );
  Span4Mux_h4 t2723 (
    .I(seg_12_12_sp4_h_l_46_35116),
    .O(seg_16_12_sp4_h_l_46_50440)
  );
  Span4Mux_h4 t2724 (
    .I(seg_8_12_sp4_h_l_46_20423),
    .O(seg_12_12_sp4_h_l_46_35116)
  );
  LocalMux t2725 (
    .I(seg_3_12_sp4_h_r_4_16595),
    .O(seg_3_12_local_g0_4_16499)
  );
  LocalMux t2726 (
    .I(seg_7_9_sp4_v_b_45_27544),
    .O(seg_7_9_local_g3_5_30848)
  );
  Span4Mux_v3 t2727 (
    .I(seg_7_12_sp4_h_l_45_16599),
    .O(seg_7_9_sp4_v_b_45_27544)
  );
  LocalMux t2728 (
    .I(seg_3_6_sp4_v_b_34_11920),
    .O(seg_3_6_local_g3_2_15783)
  );
  Span4Mux_v2 t2729 (
    .I(seg_3_8_sp4_v_t_47_12412),
    .O(seg_3_6_sp4_v_b_34_11920)
  );
  CascadeMux t273 (
    .I(net_19629),
    .O(net_19629_cascademuxed)
  );
  Span4Mux_v4 t2730 (
    .I(seg_3_12_sp4_h_r_10_16591),
    .O(seg_3_8_sp4_v_t_47_12412)
  );
  LocalMux t2731 (
    .I(seg_0_24_sp4_h_r_35_5274),
    .O(seg_0_24_local_g2_3_5134)
  );
  Span4Mux_h2 t2732 (
    .I(seg_2_24_sp4_v_b_11_9835),
    .O(seg_0_24_sp4_h_r_35_5274)
  );
  Span4Mux_v4 t2733 (
    .I(seg_2_20_sp4_v_b_8_9246),
    .O(seg_2_24_sp4_v_b_11_9835)
  );
  Span4Mux_v4 t2734 (
    .I(seg_2_16_sp4_v_b_5_8653),
    .O(seg_2_20_sp4_v_b_8_9246)
  );
  Span4Mux_v4 t2735 (
    .I(seg_2_12_sp4_h_r_11_12761),
    .O(seg_2_16_sp4_v_b_5_8653)
  );
  LocalMux t2736 (
    .I(seg_7_9_sp4_h_r_19_27531),
    .O(seg_7_9_local_g1_3_30830)
  );
  Span4Mux_h1 t2737 (
    .I(seg_6_9_sp4_v_t_43_24024),
    .O(seg_7_9_sp4_h_r_19_27531)
  );
  LocalMux t2738 (
    .I(seg_0_6_sp4_h_r_29_1406),
    .O(seg_0_6_local_g2_5_1275)
  );
  Span4Mux_h2 t2739 (
    .I(seg_2_6_sp4_h_r_9_12031),
    .O(seg_0_6_sp4_h_r_29_1406)
  );
  CascadeMux t274 (
    .I(net_19641),
    .O(net_19641_cascademuxed)
  );
  Span4Mux_h4 t2740 (
    .I(seg_6_6_sp4_v_t_38_23650),
    .O(seg_2_6_sp4_h_r_9_12031)
  );
  Span4Mux_v4 t2741 (
    .I(seg_6_10_sp4_v_t_42_24146),
    .O(seg_6_6_sp4_v_t_38_23650)
  );
  LocalMux t2742 (
    .I(seg_14_10_sp4_h_r_10_57854),
    .O(seg_14_10_local_g0_2_57760)
  );
  Span4Mux_h0 t2743 (
    .I(seg_14_10_sp4_h_l_39_42533),
    .O(seg_14_10_sp4_h_r_10_57854)
  );
  Span4Mux_h4 t2744 (
    .I(seg_10_10_sp4_h_l_39_27629),
    .O(seg_14_10_sp4_h_l_39_42533)
  );
  Span4Mux_h4 t2745 (
    .I(seg_6_10_sp4_v_t_44_24148),
    .O(seg_10_10_sp4_h_l_39_27629)
  );
  LocalMux t2746 (
    .I(seg_4_7_sp4_r_v_b_23_19582),
    .O(seg_4_7_local_g3_7_19742)
  );
  Span4Mux_v1 t2747 (
    .I(seg_5_8_sp4_v_t_39_20066),
    .O(seg_4_7_sp4_r_v_b_23_19582)
  );
  LocalMux t2748 (
    .I(seg_5_10_sp4_v_b_26_20066),
    .O(seg_5_10_local_g2_2_23929)
  );
  LocalMux t2749 (
    .I(seg_0_7_sp4_r_v_b_42_1646),
    .O(seg_0_7_local_g3_2_1486)
  );
  CascadeMux t275 (
    .I(net_19647),
    .O(net_19647_cascademuxed)
  );
  Span4Mux_v3 t2750 (
    .I(seg_1_10_sp4_h_r_2_8200),
    .O(seg_0_7_sp4_r_v_b_42_1646)
  );
  Span4Mux_h4 t2751 (
    .I(seg_5_10_sp4_v_t_39_20312),
    .O(seg_1_10_sp4_h_r_2_8200)
  );
  LocalMux t2752 (
    .I(seg_0_17_sp4_r_v_b_18_3352),
    .O(seg_0_17_local_g3_2_3606)
  );
  Span4Mux_v3 t2753 (
    .I(seg_1_14_sp4_h_r_7_8793),
    .O(seg_0_17_sp4_r_v_b_18_3352)
  );
  Span4Mux_h4 t2754 (
    .I(seg_5_14_sp4_v_b_2_20312),
    .O(seg_1_14_sp4_h_r_7_8793)
  );
  LocalMux t2755 (
    .I(seg_5_2_sp4_v_b_33_19082),
    .O(seg_5_2_local_g2_1_22944)
  );
  Span4Mux_v2 t2756 (
    .I(seg_5_4_sp4_v_t_43_19578),
    .O(seg_5_2_sp4_v_b_33_19082)
  );
  Span4Mux_v4 t2757 (
    .I(seg_5_8_sp4_v_t_43_20070),
    .O(seg_5_4_sp4_v_t_43_19578)
  );
  LocalMux t2758 (
    .I(seg_8_3_sp4_r_v_b_13_33767),
    .O(seg_8_3_local_g2_5_33933)
  );
  Span4Mux_v1 t2759 (
    .I(seg_9_4_sp4_h_l_43_23275),
    .O(seg_8_3_sp4_r_v_b_13_33767)
  );
  CascadeMux t276 (
    .I(net_19653),
    .O(net_19653_cascademuxed)
  );
  Span4Mux_h4 t2760 (
    .I(seg_5_4_sp4_v_t_43_19578),
    .O(seg_9_4_sp4_h_l_43_23275)
  );
  LocalMux t2761 (
    .I(seg_4_12_neigh_op_tnr_0_20408),
    .O(seg_4_12_local_g3_0_20350)
  );
  LocalMux t2762 (
    .I(seg_4_12_neigh_op_tnr_2_20410),
    .O(seg_4_12_local_g2_2_20344)
  );
  LocalMux t2763 (
    .I(seg_5_13_lutff_3_out_20411),
    .O(seg_5_13_local_g0_3_24283)
  );
  LocalMux t2764 (
    .I(seg_5_12_neigh_op_top_4_20412),
    .O(seg_5_12_local_g0_4_24161)
  );
  LocalMux t2765 (
    .I(seg_5_13_lutff_5_out_20413),
    .O(seg_5_13_local_g1_5_24293)
  );
  LocalMux t2766 (
    .I(seg_5_13_lutff_6_out_20414),
    .O(seg_5_13_local_g0_6_24286)
  );
  LocalMux t2767 (
    .I(seg_5_12_neigh_op_top_7_20415),
    .O(seg_5_12_local_g0_7_24164)
  );
  LocalMux t2768 (
    .I(seg_5_3_sp12_v_b_20_22861),
    .O(seg_5_3_local_g3_4_23078)
  );
  LocalMux t2769 (
    .I(seg_3_8_sp4_r_v_b_18_15869),
    .O(seg_3_8_local_g3_2_16029)
  );
  CascadeMux t277 (
    .I(net_19659),
    .O(net_19659_cascademuxed)
  );
  Span4Mux_v1 t2770 (
    .I(seg_4_9_sp4_v_t_42_16361),
    .O(seg_3_8_sp4_r_v_b_18_15869)
  );
  Span4Mux_v4 t2771 (
    .I(seg_4_13_sp4_h_r_7_20552),
    .O(seg_4_9_sp4_v_t_42_16361)
  );
  LocalMux t2772 (
    .I(seg_14_10_sp4_h_r_7_57861),
    .O(seg_14_10_local_g1_7_57773)
  );
  Span4Mux_h0 t2773 (
    .I(seg_14_10_sp4_h_l_42_42538),
    .O(seg_14_10_sp4_h_r_7_57861)
  );
  Span4Mux_h4 t2774 (
    .I(seg_10_10_sp4_h_l_41_27631),
    .O(seg_14_10_sp4_h_l_42_42538)
  );
  Span4Mux_h4 t2775 (
    .I(seg_6_10_sp4_v_t_41_24145),
    .O(seg_10_10_sp4_h_l_41_27631)
  );
  LocalMux t2776 (
    .I(seg_3_6_sp4_h_r_21_12030),
    .O(seg_3_6_local_g0_5_15762)
  );
  Span4Mux_h3 t2777 (
    .I(seg_6_6_sp4_v_t_39_23651),
    .O(seg_3_6_sp4_h_r_21_12030)
  );
  Span4Mux_v4 t2778 (
    .I(seg_6_10_sp4_v_t_43_24147),
    .O(seg_6_6_sp4_v_t_39_23651)
  );
  LocalMux t2779 (
    .I(seg_4_6_sp4_h_r_32_12030),
    .O(seg_4_6_local_g2_0_19604)
  );
  CascadeMux t278 (
    .I(net_19746),
    .O(net_19746_cascademuxed)
  );
  Span4Mux_h2 t2780 (
    .I(seg_6_6_sp4_v_t_39_23651),
    .O(seg_4_6_sp4_h_r_32_12030)
  );
  LocalMux t2781 (
    .I(seg_16_10_sp4_h_r_26_57856),
    .O(seg_16_10_local_g3_2_65445)
  );
  Span4Mux_h2 t2782 (
    .I(seg_14_10_sp4_h_l_43_42537),
    .O(seg_16_10_sp4_h_r_26_57856)
  );
  Span4Mux_h4 t2783 (
    .I(seg_10_10_sp4_h_l_43_27633),
    .O(seg_14_10_sp4_h_l_43_42537)
  );
  Span4Mux_h4 t2784 (
    .I(seg_6_10_sp4_v_t_43_24147),
    .O(seg_10_10_sp4_h_l_43_27633)
  );
  LocalMux t2785 (
    .I(seg_4_7_sp4_r_v_b_36_19817),
    .O(seg_4_7_local_g2_4_19731)
  );
  Span4Mux_v3 t2786 (
    .I(seg_5_10_sp4_v_t_40_20313),
    .O(seg_4_7_sp4_r_v_b_36_19817)
  );
  LocalMux t2787 (
    .I(seg_5_10_sp4_h_r_5_24012),
    .O(seg_5_10_local_g0_5_23916)
  );
  Span4Mux_h0 t2788 (
    .I(seg_5_10_sp4_v_t_40_20313),
    .O(seg_5_10_sp4_h_r_5_24012)
  );
  LocalMux t2789 (
    .I(seg_3_6_sp4_h_r_35_7611),
    .O(seg_3_6_local_g3_3_15784)
  );
  CascadeMux t279 (
    .I(net_19758),
    .O(net_19758_cascademuxed)
  );
  Span4Mux_h2 t2790 (
    .I(seg_5_6_sp4_v_t_40_19821),
    .O(seg_3_6_sp4_h_r_35_7611)
  );
  Span4Mux_v4 t2791 (
    .I(seg_5_10_sp4_v_t_44_20317),
    .O(seg_5_6_sp4_v_t_40_19821)
  );
  LocalMux t2792 (
    .I(seg_4_7_sp4_r_v_b_37_19818),
    .O(seg_4_7_local_g2_5_19732)
  );
  Span4Mux_v3 t2793 (
    .I(seg_5_10_sp4_v_t_44_20317),
    .O(seg_4_7_sp4_r_v_b_37_19818)
  );
  LocalMux t2794 (
    .I(seg_5_10_sp4_h_r_9_24016),
    .O(seg_5_10_local_g1_1_23920)
  );
  Span4Mux_h0 t2795 (
    .I(seg_5_10_sp4_v_t_44_20317),
    .O(seg_5_10_sp4_h_r_9_24016)
  );
  LocalMux t2796 (
    .I(seg_14_10_sp4_h_r_13_54022),
    .O(seg_14_10_local_g1_5_57771)
  );
  Span4Mux_h1 t2797 (
    .I(seg_13_10_sp4_h_l_44_38709),
    .O(seg_14_10_sp4_h_r_13_54022)
  );
  Span4Mux_h4 t2798 (
    .I(seg_9_10_sp4_h_l_44_24016),
    .O(seg_13_10_sp4_h_l_44_38709)
  );
  Span4Mux_h4 t2799 (
    .I(seg_5_10_sp4_v_t_44_20317),
    .O(seg_9_10_sp4_h_l_44_24016)
  );
  CascadeMux t28 (
    .I(net_7549),
    .O(net_7549_cascademuxed)
  );
  CascadeMux t280 (
    .I(net_19764),
    .O(net_19764_cascademuxed)
  );
  LocalMux t2800 (
    .I(seg_5_18_sp4_v_b_12_20924),
    .O(seg_5_18_local_g0_4_24899)
  );
  Span4Mux_v3 t2801 (
    .I(seg_5_15_sp4_v_b_10_20443),
    .O(seg_5_18_sp4_v_b_12_20924)
  );
  LocalMux t2802 (
    .I(seg_5_14_lutff_1_out_20532),
    .O(seg_5_14_local_g3_1_24428)
  );
  LocalMux t2803 (
    .I(seg_5_14_lutff_2_out_20533),
    .O(seg_5_14_local_g2_2_24421)
  );
  LocalMux t2804 (
    .I(seg_5_14_lutff_4_out_20535),
    .O(seg_5_14_local_g2_4_24423)
  );
  LocalMux t2805 (
    .I(seg_5_14_lutff_5_out_20536),
    .O(seg_5_14_local_g3_5_24432)
  );
  LocalMux t2806 (
    .I(seg_6_9_sp4_v_b_28_23776),
    .O(seg_6_9_local_g3_4_27477)
  );
  Span4Mux_v2 t2807 (
    .I(seg_6_11_sp4_v_t_41_24268),
    .O(seg_6_9_sp4_v_b_28_23776)
  );
  LocalMux t2808 (
    .I(seg_6_11_sp4_h_r_4_27733),
    .O(seg_6_11_local_g1_4_27665)
  );
  Span4Mux_h0 t2809 (
    .I(seg_6_11_sp4_v_t_41_24268),
    .O(seg_6_11_sp4_h_r_4_27733)
  );
  CascadeMux t281 (
    .I(net_19770),
    .O(net_19770_cascademuxed)
  );
  LocalMux t2810 (
    .I(seg_6_9_sp4_v_b_38_23896),
    .O(seg_6_9_local_g2_6_27471)
  );
  Span4Mux_v3 t2811 (
    .I(seg_6_12_sp4_v_t_42_24392),
    .O(seg_6_9_sp4_v_b_38_23896)
  );
  LocalMux t2812 (
    .I(seg_6_11_sp4_v_b_14_23896),
    .O(seg_6_11_local_g0_6_27659)
  );
  Span4Mux_v1 t2813 (
    .I(seg_6_12_sp4_v_t_42_24392),
    .O(seg_6_11_sp4_v_b_14_23896)
  );
  LocalMux t2814 (
    .I(seg_5_15_lutff_1_out_20655),
    .O(seg_5_15_local_g3_1_24551)
  );
  LocalMux t2815 (
    .I(seg_5_15_lutff_3_out_20657),
    .O(seg_5_15_local_g3_3_24553)
  );
  LocalMux t2816 (
    .I(seg_4_15_neigh_op_rgt_4_20658),
    .O(seg_4_15_local_g2_4_20715)
  );
  LocalMux t2817 (
    .I(seg_5_15_lutff_6_out_20660),
    .O(seg_5_15_local_g2_6_24548)
  );
  LocalMux t2818 (
    .I(seg_5_15_lutff_7_out_20661),
    .O(seg_5_15_local_g3_7_24557)
  );
  LocalMux t2819 (
    .I(seg_7_14_sp4_h_r_19_28041),
    .O(seg_7_14_local_g1_3_31445)
  );
  CascadeMux t282 (
    .I(net_19788),
    .O(net_19788_cascademuxed)
  );
  Span4Mux_h1 t2820 (
    .I(seg_6_14_sp4_v_t_43_24639),
    .O(seg_7_14_sp4_h_r_19_28041)
  );
  LocalMux t2821 (
    .I(seg_5_12_sp4_v_b_41_20437),
    .O(seg_5_12_local_g3_1_24182)
  );
  LocalMux t2822 (
    .I(seg_5_4_sp4_r_v_b_17_23038),
    .O(seg_5_4_local_g3_1_23198)
  );
  Span4Mux_v1 t2823 (
    .I(seg_6_5_sp4_v_t_36_23525),
    .O(seg_5_4_sp4_r_v_b_17_23038)
  );
  Span4Mux_v4 t2824 (
    .I(seg_6_9_sp4_v_t_40_24021),
    .O(seg_6_5_sp4_v_t_36_23525)
  );
  Span4Mux_v4 t2825 (
    .I(seg_6_13_sp4_v_t_39_24512),
    .O(seg_6_9_sp4_v_t_40_24021)
  );
  LocalMux t2826 (
    .I(seg_5_8_sp4_h_r_3_23764),
    .O(seg_5_8_local_g0_3_23668)
  );
  Span4Mux_h0 t2827 (
    .I(seg_5_8_sp4_v_t_47_20074),
    .O(seg_5_8_sp4_h_r_3_23764)
  );
  Span4Mux_v4 t2828 (
    .I(seg_5_12_sp4_v_t_47_20566),
    .O(seg_5_8_sp4_v_t_47_20074)
  );
  LocalMux t2829 (
    .I(seg_4_6_sp4_r_v_b_6_19332),
    .O(seg_4_6_local_g1_6_19602)
  );
  CascadeMux t283 (
    .I(net_19869),
    .O(net_19869_cascademuxed)
  );
  Span4Mux_v1 t2830 (
    .I(seg_5_6_sp4_v_t_38_19819),
    .O(seg_4_6_sp4_r_v_b_6_19332)
  );
  Span4Mux_v4 t2831 (
    .I(seg_5_10_sp4_v_t_37_20310),
    .O(seg_5_6_sp4_v_t_38_19819)
  );
  Span4Mux_v4 t2832 (
    .I(seg_5_14_sp4_v_t_41_20806),
    .O(seg_5_10_sp4_v_t_37_20310)
  );
  LocalMux t2833 (
    .I(seg_4_6_sp4_r_v_b_32_19580),
    .O(seg_4_6_local_g0_3_19591)
  );
  Span4Mux_v2 t2834 (
    .I(seg_5_8_sp4_v_t_37_20064),
    .O(seg_4_6_sp4_r_v_b_32_19580)
  );
  Span4Mux_v4 t2835 (
    .I(seg_5_12_sp4_v_t_41_20560),
    .O(seg_5_8_sp4_v_t_37_20064)
  );
  LocalMux t2836 (
    .I(seg_5_17_lutff_1_out_20901),
    .O(seg_5_17_local_g0_1_24773)
  );
  LocalMux t2837 (
    .I(seg_12_1_sp4_h_r_42_37564),
    .O(seg_12_1_local_g2_2_48968)
  );
  Span4Mux_h3 t2838 (
    .I(seg_9_1_sp4_v_t_39_33898),
    .O(seg_12_1_sp4_h_r_42_37564)
  );
  Span4Mux_v4 t2839 (
    .I(seg_9_5_sp4_v_t_43_34394),
    .O(seg_9_1_sp4_v_t_39_33898)
  );
  CascadeMux t284 (
    .I(net_19875),
    .O(net_19875_cascademuxed)
  );
  Span4Mux_v4 t2840 (
    .I(seg_9_9_sp4_v_t_47_34890),
    .O(seg_9_5_sp4_v_t_43_34394)
  );
  Span4Mux_v4 t2841 (
    .I(seg_9_13_sp4_v_t_39_35374),
    .O(seg_9_9_sp4_v_t_47_34890)
  );
  Span4Mux_v4 t2842 (
    .I(seg_9_17_sp4_h_l_39_24870),
    .O(seg_9_13_sp4_v_t_39_35374)
  );
  LocalMux t2843 (
    .I(seg_17_7_sp4_v_b_34_65044),
    .O(seg_17_7_local_g2_2_68899)
  );
  Span4Mux_v2 t2844 (
    .I(seg_17_9_sp4_h_l_47_53901),
    .O(seg_17_7_sp4_v_b_34_65044)
  );
  Span4Mux_h4 t2845 (
    .I(seg_13_9_sp4_h_l_47_38577),
    .O(seg_17_9_sp4_h_l_47_53901)
  );
  Span4Mux_h4 t2846 (
    .I(seg_9_9_sp4_v_t_47_34890),
    .O(seg_13_9_sp4_h_l_47_38577)
  );
  LocalMux t2847 (
    .I(seg_3_4_sp4_v_b_19_11547),
    .O(seg_3_4_local_g1_3_15522)
  );
  Span4Mux_v1 t2848 (
    .I(seg_3_5_sp4_v_t_43_12039),
    .O(seg_3_4_sp4_v_b_19_11547)
  );
  Span4Mux_v4 t2849 (
    .I(seg_3_9_sp4_v_t_43_12531),
    .O(seg_3_5_sp4_v_t_43_12039)
  );
  CascadeMux t285 (
    .I(net_19881),
    .O(net_19881_cascademuxed)
  );
  Span4Mux_v4 t2850 (
    .I(seg_3_13_sp4_v_t_38_13018),
    .O(seg_3_9_sp4_v_t_43_12531)
  );
  Span4Mux_v4 t2851 (
    .I(seg_3_17_sp4_h_r_10_17206),
    .O(seg_3_13_sp4_v_t_38_13018)
  );
  LocalMux t2852 (
    .I(seg_3_5_sp4_h_r_6_15736),
    .O(seg_3_5_local_g1_6_15648)
  );
  Span4Mux_h0 t2853 (
    .I(seg_3_5_sp4_v_t_43_12039),
    .O(seg_3_5_sp4_h_r_6_15736)
  );
  LocalMux t2854 (
    .I(seg_3_6_sp4_v_b_43_12039),
    .O(seg_3_6_local_g2_3_15776)
  );
  Span4Mux_v3 t2855 (
    .I(seg_3_9_sp4_v_t_43_12531),
    .O(seg_3_6_sp4_v_b_43_12039)
  );
  LocalMux t2856 (
    .I(seg_7_17_sp4_r_v_b_22_31673),
    .O(seg_7_17_local_g3_6_31833)
  );
  Span4Mux_v1 t2857 (
    .I(seg_8_18_sp4_h_l_46_21161),
    .O(seg_7_17_sp4_r_v_b_22_31673)
  );
  LocalMux t2858 (
    .I(seg_7_17_sp4_v_b_13_28148),
    .O(seg_7_17_local_g0_5_31808)
  );
  Span4Mux_v1 t2859 (
    .I(seg_7_18_sp4_h_l_37_17327),
    .O(seg_7_17_sp4_v_b_13_28148)
  );
  CascadeMux t286 (
    .I(net_19887),
    .O(net_19887_cascademuxed)
  );
  LocalMux t2860 (
    .I(seg_5_16_sp4_r_v_b_27_24634),
    .O(seg_5_16_local_g1_3_24660)
  );
  LocalMux t2861 (
    .I(seg_5_18_neigh_op_top_0_21146),
    .O(seg_5_18_local_g0_0_24895)
  );
  LocalMux t2862 (
    .I(seg_7_16_sp4_v_b_43_28256),
    .O(seg_7_16_local_g2_3_31699)
  );
  Span4Mux_v3 t2863 (
    .I(seg_7_19_sp4_h_l_37_17450),
    .O(seg_7_16_sp4_v_b_43_28256)
  );
  LocalMux t2864 (
    .I(seg_3_1_sp4_h_r_28_6843),
    .O(seg_3_1_local_g2_4_15122)
  );
  Span4Mux_h2 t2865 (
    .I(seg_5_1_sp4_v_t_47_19213),
    .O(seg_3_1_sp4_h_r_28_6843)
  );
  Span4Mux_v4 t2866 (
    .I(seg_5_5_sp4_v_t_47_19705),
    .O(seg_5_1_sp4_v_t_47_19213)
  );
  Sp12to4 t2867 (
    .I(seg_5_8_sp12_v_b_23_23635),
    .O(seg_5_5_sp4_v_t_47_19705)
  );
  Span12Mux_v11 t2868 (
    .I(seg_5_19_sp12_v_t_23_25111),
    .O(seg_5_8_sp12_v_b_23_23635)
  );
  LocalMux t2869 (
    .I(seg_3_3_sp4_h_r_26_7171),
    .O(seg_3_3_local_g3_2_15414)
  );
  CascadeMux t287 (
    .I(net_19893),
    .O(net_19893_cascademuxed)
  );
  Span4Mux_h2 t2870 (
    .I(seg_5_3_sp4_v_t_45_19457),
    .O(seg_3_3_sp4_h_r_26_7171)
  );
  Span4Mux_v4 t2871 (
    .I(seg_5_7_sp4_v_t_45_19949),
    .O(seg_5_3_sp4_v_t_45_19457)
  );
  Sp12to4 t2872 (
    .I(seg_5_10_sp12_v_b_19_23635),
    .O(seg_5_7_sp4_v_t_45_19949)
  );
  Span12Mux_v9 t2873 (
    .I(seg_5_19_sp12_v_t_23_25111),
    .O(seg_5_10_sp12_v_b_19_23635)
  );
  LocalMux t2874 (
    .I(seg_3_3_sp4_h_r_29_7174),
    .O(seg_3_3_local_g3_5_15417)
  );
  Span4Mux_h2 t2875 (
    .I(seg_5_3_sp4_v_t_46_19458),
    .O(seg_3_3_sp4_h_r_29_7174)
  );
  Span4Mux_v4 t2876 (
    .I(seg_5_7_sp4_v_t_45_19949),
    .O(seg_5_3_sp4_v_t_46_19458)
  );
  LocalMux t2877 (
    .I(seg_4_1_sp4_r_v_b_1_19044),
    .O(seg_4_1_local_g1_1_18942)
  );
  Span4Mux_v1 t2878 (
    .I(seg_5_1_sp4_v_t_47_19213),
    .O(seg_4_1_sp4_r_v_b_1_19044)
  );
  LocalMux t2879 (
    .I(seg_4_3_sp4_r_v_b_4_19064),
    .O(seg_4_3_local_g1_4_19231)
  );
  CascadeMux t288 (
    .I(net_19899),
    .O(net_19899_cascademuxed)
  );
  Sp12to4 t2880 (
    .I(seg_5_2_sp12_v_b_11_22734),
    .O(seg_4_3_sp4_r_v_b_4_19064)
  );
  Span12Mux_v5 t2881 (
    .I(seg_5_7_sp12_v_t_23_23635),
    .O(seg_5_2_sp12_v_b_11_22734)
  );
  Span12Mux_v12 t2882 (
    .I(seg_5_19_sp12_v_t_23_25111),
    .O(seg_5_7_sp12_v_t_23_23635)
  );
  LocalMux t2883 (
    .I(seg_4_4_sp4_r_v_b_23_19213),
    .O(seg_4_4_local_g3_7_19373)
  );
  Span4Mux_v1 t2884 (
    .I(seg_5_5_sp4_v_t_47_19705),
    .O(seg_4_4_sp4_r_v_b_23_19213)
  );
  LocalMux t2885 (
    .I(seg_3_2_sp4_h_r_25_7021),
    .O(seg_3_2_local_g3_1_15290)
  );
  Span4Mux_h2 t2886 (
    .I(seg_5_2_sp4_v_t_36_19325),
    .O(seg_3_2_sp4_h_r_25_7021)
  );
  Span4Mux_v4 t2887 (
    .I(seg_5_6_sp4_v_t_47_19828),
    .O(seg_5_2_sp4_v_t_36_19325)
  );
  Span4Mux_v4 t2888 (
    .I(seg_5_10_sp4_v_t_42_20315),
    .O(seg_5_6_sp4_v_t_47_19828)
  );
  Span4Mux_v4 t2889 (
    .I(seg_5_14_sp4_v_t_42_20807),
    .O(seg_5_10_sp4_v_t_42_20315)
  );
  CascadeMux t289 (
    .I(net_19905),
    .O(net_19905_cascademuxed)
  );
  Span4Mux_v4 t2890 (
    .I(seg_5_18_sp4_v_t_42_21299),
    .O(seg_5_14_sp4_v_t_42_20807)
  );
  Span4Mux_v4 t2891 (
    .I(seg_5_22_sp4_v_t_41_21790),
    .O(seg_5_18_sp4_v_t_42_21299)
  );
  Span4Mux_v4 t2892 (
    .I(seg_5_26_sp4_v_t_36_22277),
    .O(seg_5_22_sp4_v_t_41_21790)
  );
  Span4Mux_v4 t2893 (
    .I(seg_5_30_sp4_v_t_40_26489),
    .O(seg_5_26_sp4_v_t_36_22277)
  );
  LocalMux t2894 (
    .I(seg_4_3_sp4_r_v_b_13_19074),
    .O(seg_4_3_local_g2_5_19240)
  );
  IoSpan4Mux t2895 (
    .I(seg_5_0_span4_horz_r_2_22756),
    .O(seg_4_3_sp4_r_v_b_13_19074)
  );
  LocalMux t2896 (
    .I(seg_4_2_sp4_v_b_12_15230),
    .O(seg_4_2_local_g0_4_19100)
  );
  IoSpan4Mux t2897 (
    .I(seg_4_0_span4_horz_r_0_18923),
    .O(seg_4_2_sp4_v_b_12_15230)
  );
  LocalMux t2898 (
    .I(seg_3_1_sp4_h_r_16_11376),
    .O(seg_3_1_local_g1_0_15110)
  );
  Span4Mux_h3 t2899 (
    .I(seg_6_1_sp4_v_b_0_22874),
    .O(seg_3_1_sp4_h_r_16_11376)
  );
  CascadeMux t29 (
    .I(net_7561),
    .O(net_7561_cascademuxed)
  );
  CascadeMux t290 (
    .I(net_19911),
    .O(net_19911_cascademuxed)
  );
  LocalMux t2900 (
    .I(seg_3_3_sp4_h_r_20_11662),
    .O(seg_3_3_local_g0_4_15392)
  );
  Span4Mux_h3 t2901 (
    .I(seg_6_3_sp4_v_b_4_22895),
    .O(seg_3_3_sp4_h_r_20_11662)
  );
  LocalMux t2902 (
    .I(seg_5_4_neigh_op_bnr_5_23014),
    .O(seg_5_4_local_g1_5_23186)
  );
  LocalMux t2903 (
    .I(seg_5_4_neigh_op_bnr_4_23013),
    .O(seg_5_4_local_g0_4_23177)
  );
  LocalMux t2904 (
    .I(seg_5_4_neigh_op_bnr_7_23016),
    .O(seg_5_4_local_g1_7_23188)
  );
  LocalMux t2905 (
    .I(seg_5_4_neigh_op_bnr_6_23015),
    .O(seg_5_4_local_g0_6_23179)
  );
  LocalMux t2906 (
    .I(seg_5_4_neigh_op_rgt_1_23133),
    .O(seg_5_4_local_g2_1_23190)
  );
  LocalMux t2907 (
    .I(seg_5_4_neigh_op_rgt_0_23132),
    .O(seg_5_4_local_g2_0_23189)
  );
  LocalMux t2908 (
    .I(seg_3_7_sp4_v_b_12_11909),
    .O(seg_3_7_local_g0_4_15884)
  );
  Span4Mux_v3 t2909 (
    .I(seg_3_4_sp4_h_r_1_15606),
    .O(seg_3_7_sp4_v_b_12_11909)
  );
  CascadeMux t291 (
    .I(net_19992),
    .O(net_19992_cascademuxed)
  );
  LocalMux t2910 (
    .I(seg_3_7_sp4_v_b_16_11913),
    .O(seg_3_7_local_g1_0_15888)
  );
  Span4Mux_v3 t2911 (
    .I(seg_3_4_sp4_h_r_11_15608),
    .O(seg_3_7_sp4_v_b_16_11913)
  );
  LocalMux t2912 (
    .I(seg_3_7_sp4_h_r_2_15978),
    .O(seg_3_7_local_g0_2_15882)
  );
  Span4Mux_h4 t2913 (
    .I(seg_7_7_sp4_v_b_2_27028),
    .O(seg_3_7_sp4_h_r_2_15978)
  );
  LocalMux t2914 (
    .I(seg_3_7_sp4_h_r_6_15982),
    .O(seg_3_7_local_g1_6_15894)
  );
  Span4Mux_h4 t2915 (
    .I(seg_7_7_sp4_v_b_6_27032),
    .O(seg_3_7_sp4_h_r_6_15982)
  );
  LocalMux t2916 (
    .I(seg_3_7_sp4_h_r_23_12145),
    .O(seg_3_7_local_g1_7_15895)
  );
  Span4Mux_h3 t2917 (
    .I(seg_6_7_sp4_v_b_5_23283),
    .O(seg_3_7_sp4_h_r_23_12145)
  );
  LocalMux t2918 (
    .I(seg_3_7_sp4_h_r_20_12154),
    .O(seg_3_7_local_g1_4_15892)
  );
  Span4Mux_h3 t2919 (
    .I(seg_6_7_sp4_v_b_9_23287),
    .O(seg_3_7_sp4_h_r_20_12154)
  );
  CascadeMux t292 (
    .I(net_19998),
    .O(net_19998_cascademuxed)
  );
  LocalMux t2920 (
    .I(seg_5_9_neigh_op_rgt_5_23752),
    .O(seg_5_9_local_g3_5_23817)
  );
  LocalMux t2921 (
    .I(seg_5_9_neigh_op_rgt_2_23749),
    .O(seg_5_9_local_g2_2_23806)
  );
  LocalMux t2922 (
    .I(seg_5_9_neigh_op_rgt_0_23747),
    .O(seg_5_9_local_g2_0_23804)
  );
  LocalMux t2923 (
    .I(seg_1_9_sp12_h_r_5_2002),
    .O(seg_1_9_local_g1_5_7944)
  );
  LocalMux t2924 (
    .I(seg_2_9_sp12_h_r_12_2012),
    .O(seg_2_9_local_g0_4_12299)
  );
  LocalMux t2925 (
    .I(seg_1_9_sp12_h_r_13_1992),
    .O(seg_1_9_local_g0_5_7936)
  );
  LocalMux t2926 (
    .I(seg_1_9_sp4_h_r_25_2032),
    .O(seg_1_9_local_g3_1_7956)
  );
  Span4Mux_h2 t2927 (
    .I(seg_3_9_sp4_h_r_5_16227),
    .O(seg_1_9_sp4_h_r_25_2032)
  );
  LocalMux t2928 (
    .I(seg_5_11_sp4_r_v_b_10_23782),
    .O(seg_5_11_local_g2_2_24052)
  );
  LocalMux t2929 (
    .I(seg_5_9_neigh_op_tnr_7_23877),
    .O(seg_5_9_local_g2_7_23811)
  );
  CascadeMux t293 (
    .I(net_20004),
    .O(net_20004_cascademuxed)
  );
  LocalMux t2930 (
    .I(seg_5_9_neigh_op_tnr_3_23873),
    .O(seg_5_9_local_g2_3_23807)
  );
  LocalMux t2931 (
    .I(seg_5_9_neigh_op_tnr_2_23872),
    .O(seg_5_9_local_g3_2_23814)
  );
  LocalMux t2932 (
    .I(seg_5_9_neigh_op_tnr_1_23871),
    .O(seg_5_9_local_g2_1_23805)
  );
  LocalMux t2933 (
    .I(seg_5_9_neigh_op_tnr_0_23870),
    .O(seg_5_9_local_g3_0_23812)
  );
  LocalMux t2934 (
    .I(seg_1_9_sp4_r_v_b_23_7778),
    .O(seg_1_9_local_g3_7_7962)
  );
  Span4Mux_v1 t2935 (
    .I(seg_2_10_sp4_h_r_10_12514),
    .O(seg_1_9_sp4_r_v_b_23_7778)
  );
  Span4Mux_h4 t2936 (
    .I(seg_6_10_sp4_h_r_10_27627),
    .O(seg_2_10_sp4_h_r_10_12514)
  );
  LocalMux t2937 (
    .I(seg_1_9_sp4_v_b_15_1643),
    .O(seg_1_9_local_g1_7_7946)
  );
  Span4Mux_v1 t2938 (
    .I(seg_1_10_sp4_h_r_9_8207),
    .O(seg_1_9_sp4_v_b_15_1643)
  );
  Span4Mux_h4 t2939 (
    .I(seg_5_10_sp4_h_r_1_24006),
    .O(seg_1_10_sp4_h_r_9_8207)
  );
  CascadeMux t294 (
    .I(net_20010),
    .O(net_20010_cascademuxed)
  );
  LocalMux t2940 (
    .I(seg_1_9_sp4_r_v_b_22_7777),
    .O(seg_1_9_local_g3_6_7961)
  );
  Span4Mux_v1 t2941 (
    .I(seg_2_10_sp4_h_r_11_12515),
    .O(seg_1_9_sp4_r_v_b_22_7777)
  );
  Span4Mux_h4 t2942 (
    .I(seg_6_10_sp4_h_r_8_27635),
    .O(seg_2_10_sp4_h_r_11_12515)
  );
  LocalMux t2943 (
    .I(seg_5_12_neigh_op_bnr_5_23998),
    .O(seg_5_12_local_g1_5_24170)
  );
  LocalMux t2944 (
    .I(seg_5_11_neigh_op_rgt_4_23997),
    .O(seg_5_11_local_g2_4_24054)
  );
  LocalMux t2945 (
    .I(seg_5_11_neigh_op_rgt_2_23995),
    .O(seg_5_11_local_g3_2_24060)
  );
  LocalMux t2946 (
    .I(seg_5_11_neigh_op_rgt_0_23993),
    .O(seg_5_11_local_g3_0_24058)
  );
  LocalMux t2947 (
    .I(seg_3_11_sp4_h_r_15_12639),
    .O(seg_3_11_local_g1_7_16387)
  );
  Span4Mux_h3 t2948 (
    .I(seg_6_11_sp4_h_r_2_27731),
    .O(seg_3_11_sp4_h_r_15_12639)
  );
  LocalMux t2949 (
    .I(seg_3_11_sp4_h_r_3_16471),
    .O(seg_3_11_local_g0_3_16375)
  );
  CascadeMux t295 (
    .I(net_20016),
    .O(net_20016_cascademuxed)
  );
  LocalMux t2950 (
    .I(seg_4_11_sp4_h_r_20_16477),
    .O(seg_4_11_local_g1_4_20215)
  );
  LocalMux t2951 (
    .I(seg_3_11_sp4_h_r_11_16469),
    .O(seg_3_11_local_g1_3_16383)
  );
  LocalMux t2952 (
    .I(seg_5_11_neigh_op_tnr_4_24120),
    .O(seg_5_11_local_g3_4_24062)
  );
  LocalMux t2953 (
    .I(seg_5_11_neigh_op_tnr_0_24116),
    .O(seg_5_11_local_g2_0_24050)
  );
  LocalMux t2954 (
    .I(seg_4_11_sp4_r_v_b_21_20072),
    .O(seg_4_11_local_g3_5_20232)
  );
  Span4Mux_v1 t2955 (
    .I(seg_5_12_sp4_h_r_3_24256),
    .O(seg_4_11_sp4_r_v_b_21_20072)
  );
  LocalMux t2956 (
    .I(seg_4_11_sp4_v_b_20_16240),
    .O(seg_4_11_local_g0_4_20207)
  );
  Span4Mux_v1 t2957 (
    .I(seg_4_12_sp4_h_r_4_20426),
    .O(seg_4_11_sp4_v_b_20_16240)
  );
  LocalMux t2958 (
    .I(seg_3_11_sp4_r_v_b_14_16234),
    .O(seg_3_11_local_g2_6_16394)
  );
  Span4Mux_v1 t2959 (
    .I(seg_4_12_sp4_h_r_10_20422),
    .O(seg_3_11_sp4_r_v_b_14_16234)
  );
  CascadeMux t296 (
    .I(net_20022),
    .O(net_20022_cascademuxed)
  );
  LocalMux t2960 (
    .I(seg_1_11_sp4_r_v_b_14_8063),
    .O(seg_1_11_local_g2_6_8247)
  );
  Span4Mux_v1 t2961 (
    .I(seg_2_12_sp4_h_r_3_12763),
    .O(seg_1_11_sp4_r_v_b_14_8063)
  );
  Span4Mux_h4 t2962 (
    .I(seg_6_12_sp4_v_b_10_23905),
    .O(seg_2_12_sp4_h_r_3_12763)
  );
  LocalMux t2963 (
    .I(seg_4_11_sp4_h_r_25_12636),
    .O(seg_4_11_local_g3_1_20228)
  );
  Span4Mux_h2 t2964 (
    .I(seg_6_11_sp4_v_t_36_24263),
    .O(seg_4_11_sp4_h_r_25_12636)
  );
  LocalMux t2965 (
    .I(seg_3_11_sp4_h_r_14_12640),
    .O(seg_3_11_local_g1_6_16386)
  );
  Span4Mux_h3 t2966 (
    .I(seg_6_11_sp4_v_t_38_24265),
    .O(seg_3_11_sp4_h_r_14_12640)
  );
  LocalMux t2967 (
    .I(seg_4_3_sp4_h_r_28_11657),
    .O(seg_4_3_local_g3_4_19247)
  );
  Span4Mux_h2 t2968 (
    .I(seg_6_3_sp4_v_t_41_23284),
    .O(seg_4_3_sp4_h_r_28_11657)
  );
  Span4Mux_v4 t2969 (
    .I(seg_6_7_sp4_v_t_45_23780),
    .O(seg_6_3_sp4_v_t_41_23284)
  );
  CascadeMux t297 (
    .I(net_20028),
    .O(net_20028_cascademuxed)
  );
  Sp12to4 t2970 (
    .I(seg_6_10_sp12_v_b_19_27318),
    .O(seg_6_7_sp4_v_t_45_23780)
  );
  Span12Mux_v9 t2971 (
    .I(seg_6_19_sp12_v_t_23_28542),
    .O(seg_6_10_sp12_v_b_19_27318)
  );
  LocalMux t2972 (
    .I(seg_4_4_sp4_h_r_29_11781),
    .O(seg_4_4_local_g3_5_19371)
  );
  Span4Mux_h2 t2973 (
    .I(seg_6_4_sp4_v_t_46_23412),
    .O(seg_4_4_sp4_h_r_29_11781)
  );
  Span4Mux_v4 t2974 (
    .I(seg_6_8_sp4_v_t_45_23903),
    .O(seg_6_4_sp4_v_t_46_23412)
  );
  Span4Mux_v4 t2975 (
    .I(seg_6_12_sp4_v_t_45_24395),
    .O(seg_6_8_sp4_v_t_45_23903)
  );
  Span4Mux_v4 t2976 (
    .I(seg_6_16_sp4_v_t_40_24882),
    .O(seg_6_12_sp4_v_t_45_24395)
  );
  Span4Mux_v4 t2977 (
    .I(seg_6_20_sp4_v_t_40_25374),
    .O(seg_6_16_sp4_v_t_40_24882)
  );
  Span4Mux_v4 t2978 (
    .I(seg_6_24_sp4_v_t_40_25866),
    .O(seg_6_20_sp4_v_t_40_25374)
  );
  Span4Mux_v4 t2979 (
    .I(seg_6_28_sp4_v_t_40_26358),
    .O(seg_6_24_sp4_v_t_40_25866)
  );
  CascadeMux t298 (
    .I(net_20034),
    .O(net_20034_cascademuxed)
  );
  LocalMux t2980 (
    .I(seg_4_2_sp4_h_r_26_11532),
    .O(seg_4_2_local_g3_2_19122)
  );
  Span4Mux_h2 t2981 (
    .I(seg_6_2_sp4_v_t_45_23165),
    .O(seg_4_2_sp4_h_r_26_11532)
  );
  Span4Mux_v4 t2982 (
    .I(seg_6_6_sp4_v_t_45_23657),
    .O(seg_6_2_sp4_v_t_45_23165)
  );
  Span4Mux_v4 t2983 (
    .I(seg_6_10_sp4_v_t_45_24149),
    .O(seg_6_6_sp4_v_t_45_23657)
  );
  Span4Mux_v4 t2984 (
    .I(seg_6_14_sp4_v_t_37_24633),
    .O(seg_6_10_sp4_v_t_45_24149)
  );
  Span4Mux_v4 t2985 (
    .I(seg_6_18_sp4_v_t_37_25125),
    .O(seg_6_14_sp4_v_t_37_24633)
  );
  Span4Mux_v4 t2986 (
    .I(seg_6_22_sp4_v_t_41_25621),
    .O(seg_6_18_sp4_v_t_37_25125)
  );
  Span4Mux_v4 t2987 (
    .I(seg_6_26_sp4_v_t_36_26108),
    .O(seg_6_22_sp4_v_t_41_25621)
  );
  Span4Mux_v4 t2988 (
    .I(seg_6_30_sp4_v_t_40_29689),
    .O(seg_6_26_sp4_v_t_36_26108)
  );
  LocalMux t2989 (
    .I(seg_8_1_neigh_op_lft_1_26554),
    .O(seg_8_1_local_g1_1_33635)
  );
  CascadeMux t299 (
    .I(net_20115),
    .O(net_20115_cascademuxed)
  );
  LocalMux t2990 (
    .I(seg_8_1_neigh_op_tnl_2_26631),
    .O(seg_8_1_local_g3_2_33652)
  );
  LocalMux t2991 (
    .I(seg_7_2_lutff_3_out_26632),
    .O(seg_7_2_local_g0_3_29961)
  );
  LocalMux t2992 (
    .I(seg_8_1_neigh_op_tnl_4_26633),
    .O(seg_8_1_local_g2_4_33646)
  );
  LocalMux t2993 (
    .I(seg_7_3_lutff_2_out_26769),
    .O(seg_7_3_local_g1_2_30091)
  );
  LocalMux t2994 (
    .I(seg_10_3_sp4_h_r_37_30175),
    .O(seg_10_3_local_g2_5_41595)
  );
  LocalMux t2995 (
    .I(seg_10_3_sp4_h_r_2_41672),
    .O(seg_10_3_local_g1_2_41584)
  );
  Span4Mux_h0 t2996 (
    .I(seg_10_3_sp4_h_l_46_26914),
    .O(seg_10_3_sp4_h_r_2_41672)
  );
  LocalMux t2997 (
    .I(seg_10_3_sp4_h_r_45_30185),
    .O(seg_10_3_local_g3_5_41603)
  );
  LocalMux t2998 (
    .I(seg_7_3_neigh_op_top_0_26869),
    .O(seg_7_3_local_g0_0_30081)
  );
  LocalMux t2999 (
    .I(seg_7_4_lutff_1_out_26870),
    .O(seg_7_4_local_g2_1_30221)
  );
  CascadeMux t30 (
    .I(net_7861),
    .O(net_7861_cascademuxed)
  );
  CascadeMux t300 (
    .I(net_20121),
    .O(net_20121_cascademuxed)
  );
  LocalMux t3000 (
    .I(seg_7_5_neigh_op_bot_2_26871),
    .O(seg_7_5_local_g1_2_30337)
  );
  LocalMux t3001 (
    .I(seg_0_12_sp4_v_b_6_1868),
    .O(seg_0_12_local_g0_6_2526)
  );
  Span4Mux_v4 t3002 (
    .I(seg_0_8_sp4_h_r_6_1845),
    .O(seg_0_12_sp4_v_b_6_1868)
  );
  Span4Mux_h4 t3003 (
    .I(seg_4_8_sp4_v_b_1_15740),
    .O(seg_0_8_sp4_h_r_6_1845)
  );
  Span4Mux_v4 t3004 (
    .I(seg_4_4_sp4_h_r_7_19445),
    .O(seg_4_8_sp4_v_b_1_15740)
  );
  LocalMux t3005 (
    .I(seg_0_25_sp4_v_b_15_4892),
    .O(seg_0_25_local_g1_7_5336)
  );
  Span4Mux_v3 t3006 (
    .I(seg_0_22_sp4_h_r_8_4875),
    .O(seg_0_25_sp4_v_b_15_4892)
  );
  Span4Mux_h4 t3007 (
    .I(seg_4_22_sp4_h_r_5_21657),
    .O(seg_0_22_sp4_h_r_8_4875)
  );
  Span4Mux_h4 t3008 (
    .I(seg_8_22_sp4_v_b_0_32156),
    .O(seg_4_22_sp4_h_r_5_21657)
  );
  Span4Mux_v4 t3009 (
    .I(seg_8_18_sp4_v_b_9_31671),
    .O(seg_8_22_sp4_v_b_0_32156)
  );
  CascadeMux t301 (
    .I(net_20127),
    .O(net_20127_cascademuxed)
  );
  Span4Mux_v4 t3010 (
    .I(seg_8_14_sp4_v_b_6_31178),
    .O(seg_8_18_sp4_v_b_9_31671)
  );
  Span4Mux_v4 t3011 (
    .I(seg_8_10_sp4_v_b_3_30681),
    .O(seg_8_14_sp4_v_b_6_31178)
  );
  Span4Mux_v4 t3012 (
    .I(seg_8_6_sp4_v_b_3_30189),
    .O(seg_8_10_sp4_v_b_3_30681)
  );
  LocalMux t3013 (
    .I(seg_10_3_sp4_h_r_27_34011),
    .O(seg_10_3_local_g2_3_41593)
  );
  Span4Mux_h2 t3014 (
    .I(seg_8_3_sp4_v_t_47_30321),
    .O(seg_10_3_sp4_h_r_27_34011)
  );
  LocalMux t3015 (
    .I(seg_7_2_sp4_v_b_30_26721),
    .O(seg_7_2_local_g2_6_29980)
  );
  LocalMux t3016 (
    .I(seg_7_6_neigh_op_bot_1_26972),
    .O(seg_7_6_local_g1_1_30459)
  );
  LocalMux t3017 (
    .I(seg_7_6_neigh_op_bot_2_26973),
    .O(seg_7_6_local_g1_2_30460)
  );
  LocalMux t3018 (
    .I(seg_7_6_neigh_op_bot_3_26974),
    .O(seg_7_6_local_g0_3_30453)
  );
  LocalMux t3019 (
    .I(seg_7_6_neigh_op_bot_5_26976),
    .O(seg_7_6_local_g1_5_30463)
  );
  CascadeMux t302 (
    .I(net_20133),
    .O(net_20133_cascademuxed)
  );
  LocalMux t3020 (
    .I(seg_7_5_lutff_7_out_26978),
    .O(seg_7_5_local_g1_7_30342)
  );
  LocalMux t3021 (
    .I(seg_5_17_sp4_v_b_3_20680),
    .O(seg_5_17_local_g1_3_24783)
  );
  Span4Mux_v4 t3022 (
    .I(seg_5_13_sp4_v_b_3_20188),
    .O(seg_5_17_sp4_v_b_3_20680)
  );
  Span4Mux_v4 t3023 (
    .I(seg_5_9_sp4_v_b_0_19695),
    .O(seg_5_13_sp4_v_b_3_20188)
  );
  Span4Mux_v4 t3024 (
    .I(seg_5_5_sp4_h_r_0_23390),
    .O(seg_5_9_sp4_v_b_0_19695)
  );
  LocalMux t3025 (
    .I(seg_16_3_sp4_h_r_2_64656),
    .O(seg_16_3_local_g0_2_64560)
  );
  Span4Mux_h0 t3026 (
    .I(seg_16_3_sp4_h_l_43_49338),
    .O(seg_16_3_sp4_h_r_2_64656)
  );
  Span4Mux_h4 t3027 (
    .I(seg_12_3_sp4_h_l_43_34014),
    .O(seg_16_3_sp4_h_l_43_49338)
  );
  Span4Mux_h4 t3028 (
    .I(seg_8_3_sp4_v_t_36_30310),
    .O(seg_12_3_sp4_h_l_43_34014)
  );
  LocalMux t3029 (
    .I(seg_7_15_sp4_v_b_13_27944),
    .O(seg_7_15_local_g1_5_31570)
  );
  CascadeMux t303 (
    .I(net_20139),
    .O(net_20139_cascademuxed)
  );
  Span4Mux_v3 t3030 (
    .I(seg_7_12_sp4_v_b_0_27536),
    .O(seg_7_15_sp4_v_b_13_27944)
  );
  Span4Mux_v4 t3031 (
    .I(seg_7_8_sp4_v_b_9_27135),
    .O(seg_7_12_sp4_v_b_0_27536)
  );
  LocalMux t3032 (
    .I(seg_7_6_lutff_2_out_27075),
    .O(seg_7_6_local_g3_2_30476)
  );
  LocalMux t3033 (
    .I(seg_7_6_lutff_3_out_27076),
    .O(seg_7_6_local_g1_3_30461)
  );
  LocalMux t3034 (
    .I(seg_7_6_lutff_7_out_27080),
    .O(seg_7_6_local_g3_7_30481)
  );
  LocalMux t3035 (
    .I(seg_0_7_sp4_r_v_b_45_1649),
    .O(seg_0_7_local_g3_5_1489)
  );
  Span4Mux_v1 t3036 (
    .I(seg_1_6_sp4_h_r_2_7612),
    .O(seg_0_7_sp4_r_v_b_45_1649)
  );
  Span4Mux_h4 t3037 (
    .I(seg_5_6_sp4_h_r_2_23517),
    .O(seg_1_6_sp4_h_r_2_7612)
  );
  LocalMux t3038 (
    .I(seg_2_6_sp4_h_r_12_7609),
    .O(seg_2_6_local_g0_4_11930)
  );
  Span4Mux_h3 t3039 (
    .I(seg_5_6_sp4_h_r_10_23515),
    .O(seg_2_6_sp4_h_r_12_7609)
  );
  CascadeMux t304 (
    .I(net_20145),
    .O(net_20145_cascademuxed)
  );
  LocalMux t3040 (
    .I(seg_0_7_sp4_v_b_40_1448),
    .O(seg_0_7_local_g3_0_1484)
  );
  Span4Mux_v1 t3041 (
    .I(seg_0_6_sp4_h_r_5_1427),
    .O(seg_0_7_sp4_v_b_40_1448)
  );
  Span4Mux_h4 t3042 (
    .I(seg_4_6_sp4_h_r_5_19689),
    .O(seg_0_6_sp4_h_r_5_1427)
  );
  LocalMux t3043 (
    .I(seg_0_17_sp4_v_b_23_3159),
    .O(seg_0_17_local_g0_7_3587)
  );
  Span4Mux_v3 t3044 (
    .I(seg_0_14_sp4_v_b_7_2304),
    .O(seg_0_17_sp4_v_b_23_3159)
  );
  Span4Mux_v4 t3045 (
    .I(seg_0_10_sp4_v_b_11_1454),
    .O(seg_0_14_sp4_v_b_7_2304)
  );
  Span4Mux_v4 t3046 (
    .I(seg_0_6_sp4_h_r_5_1427),
    .O(seg_0_10_sp4_v_b_11_1454)
  );
  LocalMux t3047 (
    .I(seg_0_17_sp4_v_b_18_3154),
    .O(seg_0_17_local_g1_2_3590)
  );
  Span4Mux_v3 t3048 (
    .I(seg_0_14_sp4_v_b_11_2308),
    .O(seg_0_17_sp4_v_b_18_3154)
  );
  Span4Mux_v4 t3049 (
    .I(seg_0_10_sp4_v_b_3_1446),
    .O(seg_0_14_sp4_v_b_11_2308)
  );
  CascadeMux t305 (
    .I(net_20151),
    .O(net_20151_cascademuxed)
  );
  Span4Mux_v4 t3050 (
    .I(seg_0_6_sp4_h_r_9_1431),
    .O(seg_0_10_sp4_v_b_3_1446)
  );
  Span4Mux_h4 t3051 (
    .I(seg_4_6_sp4_h_r_9_19693),
    .O(seg_0_6_sp4_h_r_9_1431)
  );
  LocalMux t3052 (
    .I(seg_0_7_sp4_h_r_17_1601),
    .O(seg_0_7_local_g0_1_1461)
  );
  Span4Mux_h3 t3053 (
    .I(seg_3_7_sp4_h_r_1_15975),
    .O(seg_0_7_sp4_h_r_17_1601)
  );
  Span4Mux_h4 t3054 (
    .I(seg_7_7_sp4_v_b_1_27025),
    .O(seg_3_7_sp4_h_r_1_15975)
  );
  LocalMux t3055 (
    .I(seg_0_17_sp4_h_r_18_3722),
    .O(seg_0_17_local_g0_2_3582)
  );
  Span4Mux_h3 t3056 (
    .I(seg_3_17_sp4_v_b_7_13022),
    .O(seg_0_17_sp4_h_r_18_3722)
  );
  Span4Mux_v4 t3057 (
    .I(seg_3_13_sp4_h_r_7_16721),
    .O(seg_3_17_sp4_v_b_7_13022)
  );
  Span4Mux_h4 t3058 (
    .I(seg_7_13_sp4_v_b_7_27643),
    .O(seg_3_13_sp4_h_r_7_16721)
  );
  Span4Mux_v4 t3059 (
    .I(seg_7_9_sp4_v_b_7_27235),
    .O(seg_7_13_sp4_v_b_7_27643)
  );
  CascadeMux t306 (
    .I(net_20262),
    .O(net_20262_cascademuxed)
  );
  LocalMux t3060 (
    .I(seg_7_8_neigh_op_bot_0_27175),
    .O(seg_7_8_local_g1_0_30704)
  );
  LocalMux t3061 (
    .I(seg_8_8_neigh_op_bnl_1_27176),
    .O(seg_8_8_local_g2_1_34544)
  );
  LocalMux t3062 (
    .I(seg_7_7_lutff_2_out_27177),
    .O(seg_7_7_local_g2_2_30591)
  );
  LocalMux t3063 (
    .I(seg_7_7_lutff_3_out_27178),
    .O(seg_7_7_local_g2_3_30592)
  );
  LocalMux t3064 (
    .I(seg_7_8_neigh_op_bot_6_27181),
    .O(seg_7_8_local_g0_6_30702)
  );
  LocalMux t3065 (
    .I(seg_7_7_lutff_7_out_27182),
    .O(seg_7_7_local_g0_7_30580)
  );
  LocalMux t3066 (
    .I(seg_5_6_sp4_v_b_13_19449),
    .O(seg_5_6_local_g0_5_23424)
  );
  Span4Mux_v1 t3067 (
    .I(seg_5_7_sp4_h_r_0_23636),
    .O(seg_5_6_sp4_v_b_13_19449)
  );
  LocalMux t3068 (
    .I(seg_5_6_sp4_v_b_15_19451),
    .O(seg_5_6_local_g0_7_23426)
  );
  Span4Mux_v1 t3069 (
    .I(seg_5_7_sp4_h_r_2_23640),
    .O(seg_5_6_sp4_v_b_15_19451)
  );
  CascadeMux t307 (
    .I(net_20274),
    .O(net_20274_cascademuxed)
  );
  LocalMux t3070 (
    .I(seg_7_8_lutff_0_out_27277),
    .O(seg_7_8_local_g0_0_30696)
  );
  LocalMux t3071 (
    .I(seg_8_8_neigh_op_lft_1_27278),
    .O(seg_8_8_local_g0_1_34528)
  );
  LocalMux t3072 (
    .I(seg_8_8_neigh_op_lft_2_27279),
    .O(seg_8_8_local_g0_2_34529)
  );
  LocalMux t3073 (
    .I(seg_8_8_neigh_op_lft_4_27281),
    .O(seg_8_8_local_g0_4_34531)
  );
  LocalMux t3074 (
    .I(seg_8_8_neigh_op_lft_5_27282),
    .O(seg_8_8_local_g0_5_34532)
  );
  LocalMux t3075 (
    .I(seg_8_8_neigh_op_lft_6_27283),
    .O(seg_8_8_local_g1_6_34541)
  );
  LocalMux t3076 (
    .I(seg_8_8_neigh_op_lft_7_27284),
    .O(seg_8_8_local_g0_7_34534)
  );
  LocalMux t3077 (
    .I(seg_7_11_sp4_v_b_3_27435),
    .O(seg_7_11_local_g1_3_31076)
  );
  LocalMux t3078 (
    .I(seg_7_15_sp12_v_b_2_30296),
    .O(seg_7_15_local_g3_2_31583)
  );
  LocalMux t3079 (
    .I(seg_7_15_sp12_v_b_4_30420),
    .O(seg_7_15_local_g2_4_31577)
  );
  CascadeMux t308 (
    .I(net_20367),
    .O(net_20367_cascademuxed)
  );
  LocalMux t3080 (
    .I(seg_5_16_sp4_r_v_b_18_24515),
    .O(seg_5_16_local_g3_2_24675)
  );
  Span4Mux_v3 t3081 (
    .I(seg_6_13_sp4_v_b_7_24023),
    .O(seg_5_16_sp4_r_v_b_18_24515)
  );
  Span4Mux_v4 t3082 (
    .I(seg_6_9_sp4_h_r_1_27524),
    .O(seg_6_13_sp4_v_b_7_24023)
  );
  LocalMux t3083 (
    .I(seg_5_16_sp4_v_b_20_20686),
    .O(seg_5_16_local_g0_4_24653)
  );
  Span4Mux_v3 t3084 (
    .I(seg_5_13_sp4_v_b_6_20193),
    .O(seg_5_16_sp4_v_b_20_20686)
  );
  Span4Mux_v4 t3085 (
    .I(seg_5_9_sp4_h_r_0_23882),
    .O(seg_5_13_sp4_v_b_6_20193)
  );
  LocalMux t3086 (
    .I(seg_7_15_sp4_v_b_1_27841),
    .O(seg_7_15_local_g0_1_31558)
  );
  Span4Mux_v4 t3087 (
    .I(seg_7_11_sp4_v_b_10_27444),
    .O(seg_7_15_sp4_v_b_1_27841)
  );
  LocalMux t3088 (
    .I(seg_7_15_sp4_v_b_17_27948),
    .O(seg_7_15_local_g1_1_31566)
  );
  Span4Mux_v3 t3089 (
    .I(seg_7_12_sp4_v_b_1_27535),
    .O(seg_7_15_sp4_v_b_17_27948)
  );
  CascadeMux t309 (
    .I(net_20391),
    .O(net_20391_cascademuxed)
  );
  LocalMux t3090 (
    .I(seg_7_15_sp4_v_b_14_27945),
    .O(seg_7_15_local_g0_6_31563)
  );
  Span4Mux_v3 t3091 (
    .I(seg_7_12_sp4_v_b_3_27537),
    .O(seg_7_15_sp4_v_b_14_27945)
  );
  LocalMux t3092 (
    .I(seg_7_10_lutff_0_out_27481),
    .O(seg_7_10_local_g1_0_30950)
  );
  LocalMux t3093 (
    .I(seg_7_10_lutff_1_out_27482),
    .O(seg_7_10_local_g2_1_30959)
  );
  LocalMux t3094 (
    .I(seg_8_9_neigh_op_tnl_2_27483),
    .O(seg_8_9_local_g2_2_34668)
  );
  LocalMux t3095 (
    .I(seg_8_9_neigh_op_tnl_4_27485),
    .O(seg_8_9_local_g3_4_34678)
  );
  LocalMux t3096 (
    .I(seg_7_11_neigh_op_bot_6_27487),
    .O(seg_7_11_local_g0_6_31071)
  );
  LocalMux t3097 (
    .I(seg_7_13_sp4_v_b_11_27647),
    .O(seg_7_13_local_g0_3_31314)
  );
  LocalMux t3098 (
    .I(seg_7_8_sp4_v_b_30_27338),
    .O(seg_7_8_local_g3_6_30726)
  );
  LocalMux t3099 (
    .I(seg_7_12_neigh_op_bot_0_27583),
    .O(seg_7_12_local_g1_0_31196)
  );
  CascadeMux t31 (
    .I(net_7966),
    .O(net_7966_cascademuxed)
  );
  CascadeMux t310 (
    .I(net_20484),
    .O(net_20484_cascademuxed)
  );
  LocalMux t3100 (
    .I(seg_7_12_neigh_op_bot_1_27584),
    .O(seg_7_12_local_g0_1_31189)
  );
  LocalMux t3101 (
    .I(seg_7_12_neigh_op_bot_2_27585),
    .O(seg_7_12_local_g0_2_31190)
  );
  LocalMux t3102 (
    .I(seg_7_12_neigh_op_bot_3_27586),
    .O(seg_7_12_local_g1_3_31199)
  );
  LocalMux t3103 (
    .I(seg_7_11_lutff_6_out_27589),
    .O(seg_7_11_local_g1_6_31079)
  );
  LocalMux t3104 (
    .I(seg_7_12_neigh_op_bot_7_27590),
    .O(seg_7_12_local_g1_7_31203)
  );
  LocalMux t3105 (
    .I(seg_7_13_sp4_v_b_2_27640),
    .O(seg_7_13_local_g0_2_31313)
  );
  LocalMux t3106 (
    .I(seg_7_13_sp4_v_b_16_27743),
    .O(seg_7_13_local_g1_0_31319)
  );
  LocalMux t3107 (
    .I(seg_8_12_neigh_op_lft_1_27686),
    .O(seg_8_12_local_g1_1_35028)
  );
  LocalMux t3108 (
    .I(seg_8_12_neigh_op_lft_2_27687),
    .O(seg_8_12_local_g0_2_35021)
  );
  LocalMux t3109 (
    .I(seg_8_12_neigh_op_lft_3_27688),
    .O(seg_8_12_local_g1_3_35030)
  );
  CascadeMux t311 (
    .I(net_20490),
    .O(net_20490_cascademuxed)
  );
  LocalMux t3110 (
    .I(seg_8_12_neigh_op_lft_4_27689),
    .O(seg_8_12_local_g0_4_35023)
  );
  LocalMux t3111 (
    .I(seg_8_12_neigh_op_lft_5_27690),
    .O(seg_8_12_local_g1_5_35032)
  );
  LocalMux t3112 (
    .I(seg_8_12_neigh_op_lft_6_27691),
    .O(seg_8_12_local_g1_6_35033)
  );
  LocalMux t3113 (
    .I(seg_8_12_neigh_op_lft_7_27692),
    .O(seg_8_12_local_g1_7_35034)
  );
  LocalMux t3114 (
    .I(seg_8_12_neigh_op_tnl_0_27787),
    .O(seg_8_12_local_g2_0_35035)
  );
  LocalMux t3115 (
    .I(seg_7_13_lutff_1_out_27788),
    .O(seg_7_13_local_g0_1_31312)
  );
  LocalMux t3116 (
    .I(seg_7_12_neigh_op_top_2_27789),
    .O(seg_7_12_local_g1_2_31198)
  );
  LocalMux t3117 (
    .I(seg_7_12_neigh_op_top_4_27791),
    .O(seg_7_12_local_g0_4_31192)
  );
  LocalMux t3118 (
    .I(seg_7_12_neigh_op_top_5_27792),
    .O(seg_7_12_local_g1_5_31201)
  );
  LocalMux t3119 (
    .I(seg_7_12_neigh_op_top_7_27794),
    .O(seg_7_12_local_g0_7_31195)
  );
  CascadeMux t312 (
    .I(net_20496),
    .O(net_20496_cascademuxed)
  );
  LocalMux t3120 (
    .I(seg_8_3_sp4_v_b_37_30188),
    .O(seg_8_3_local_g3_5_33941)
  );
  Span4Mux_v3 t3121 (
    .I(seg_8_6_sp4_v_t_37_30680),
    .O(seg_8_3_sp4_v_b_37_30188)
  );
  Span4Mux_v4 t3122 (
    .I(seg_8_10_sp4_v_t_37_31172),
    .O(seg_8_6_sp4_v_t_37_30680)
  );
  LocalMux t3123 (
    .I(seg_8_6_sp4_h_r_5_34382),
    .O(seg_8_6_local_g0_5_34286)
  );
  Span4Mux_h0 t3124 (
    .I(seg_8_6_sp4_v_t_37_30680),
    .O(seg_8_6_sp4_h_r_5_34382)
  );
  LocalMux t3125 (
    .I(seg_9_2_sp4_h_r_13_33883),
    .O(seg_9_2_local_g1_5_37633)
  );
  Span4Mux_h1 t3126 (
    .I(seg_8_2_sp4_v_t_37_30188),
    .O(seg_9_2_sp4_h_r_13_33883)
  );
  Span4Mux_v4 t3127 (
    .I(seg_8_6_sp4_v_t_37_30680),
    .O(seg_8_2_sp4_v_t_37_30188)
  );
  LocalMux t3128 (
    .I(seg_16_10_sp4_h_r_9_65524),
    .O(seg_16_10_local_g1_1_65428)
  );
  Span4Mux_h0 t3129 (
    .I(seg_16_10_sp4_h_l_36_50192),
    .O(seg_16_10_sp4_h_r_9_65524)
  );
  CascadeMux t313 (
    .I(net_20502),
    .O(net_20502_cascademuxed)
  );
  Span4Mux_h4 t3130 (
    .I(seg_12_10_sp4_h_l_40_34874),
    .O(seg_16_10_sp4_h_l_36_50192)
  );
  Span4Mux_h4 t3131 (
    .I(seg_8_10_sp4_v_t_37_31172),
    .O(seg_12_10_sp4_h_l_40_34874)
  );
  LocalMux t3132 (
    .I(seg_7_12_sp4_r_v_b_18_31054),
    .O(seg_7_12_local_g3_2_31214)
  );
  LocalMux t3133 (
    .I(seg_7_9_sp4_v_b_17_27336),
    .O(seg_7_9_local_g1_1_30828)
  );
  Span4Mux_v1 t3134 (
    .I(seg_7_10_sp4_v_t_36_27739),
    .O(seg_7_9_sp4_v_b_17_27336)
  );
  LocalMux t3135 (
    .I(seg_7_14_lutff_6_out_27895),
    .O(seg_7_14_local_g1_6_31448)
  );
  LocalMux t3136 (
    .I(seg_8_13_neigh_op_tnl_7_27896),
    .O(seg_8_13_local_g3_7_35173)
  );
  LocalMux t3137 (
    .I(seg_9_4_sp4_r_v_b_31_37855),
    .O(seg_9_4_local_g0_7_37873)
  );
  Span4Mux_v2 t3138 (
    .I(seg_10_6_sp4_v_t_42_38347),
    .O(seg_9_4_sp4_r_v_b_31_37855)
  );
  Span4Mux_v4 t3139 (
    .I(seg_10_10_sp4_v_t_46_38843),
    .O(seg_10_6_sp4_v_t_42_38347)
  );
  CascadeMux t314 (
    .I(net_20508),
    .O(net_20508_cascademuxed)
  );
  Span4Mux_v4 t3140 (
    .I(seg_10_14_sp4_h_l_46_28036),
    .O(seg_10_10_sp4_v_t_46_38843)
  );
  LocalMux t3141 (
    .I(seg_7_5_sp4_r_v_b_19_30194),
    .O(seg_7_5_local_g3_3_30354)
  );
  Span4Mux_v1 t3142 (
    .I(seg_8_6_sp4_v_t_47_30690),
    .O(seg_7_5_sp4_r_v_b_19_30194)
  );
  Span4Mux_v4 t3143 (
    .I(seg_8_10_sp4_v_t_42_31177),
    .O(seg_8_6_sp4_v_t_47_30690)
  );
  LocalMux t3144 (
    .I(seg_8_6_sp4_h_r_3_34380),
    .O(seg_8_6_local_g0_3_34284)
  );
  Span4Mux_h0 t3145 (
    .I(seg_8_6_sp4_v_t_47_30690),
    .O(seg_8_6_sp4_h_r_3_34380)
  );
  LocalMux t3146 (
    .I(seg_16_10_sp4_h_r_4_65519),
    .O(seg_16_10_local_g0_4_65423)
  );
  Span4Mux_h0 t3147 (
    .I(seg_16_10_sp4_h_l_45_50201),
    .O(seg_16_10_sp4_h_r_4_65519)
  );
  Span4Mux_h4 t3148 (
    .I(seg_12_10_sp4_h_l_37_34867),
    .O(seg_16_10_sp4_h_l_45_50201)
  );
  Span4Mux_h4 t3149 (
    .I(seg_8_10_sp4_v_t_42_31177),
    .O(seg_12_10_sp4_h_l_37_34867)
  );
  CascadeMux t315 (
    .I(net_20514),
    .O(net_20514_cascademuxed)
  );
  LocalMux t3150 (
    .I(seg_8_11_sp4_v_b_44_31179),
    .O(seg_8_11_local_g2_4_34916)
  );
  LocalMux t3151 (
    .I(seg_7_9_sp4_v_b_20_27339),
    .O(seg_7_9_local_g1_4_30831)
  );
  Span4Mux_v1 t3152 (
    .I(seg_7_10_sp4_v_t_43_27746),
    .O(seg_7_9_sp4_v_b_20_27339)
  );
  LocalMux t3153 (
    .I(seg_7_14_neigh_op_top_2_27993),
    .O(seg_7_14_local_g1_2_31444)
  );
  LocalMux t3154 (
    .I(seg_8_5_sp4_v_b_31_30316),
    .O(seg_8_5_local_g3_7_34189)
  );
  Span4Mux_v2 t3155 (
    .I(seg_8_7_sp4_v_t_42_30808),
    .O(seg_8_5_sp4_v_b_31_30316)
  );
  Span4Mux_v4 t3156 (
    .I(seg_8_11_sp4_v_t_46_31304),
    .O(seg_8_7_sp4_v_t_42_30808)
  );
  LocalMux t3157 (
    .I(seg_9_5_sp4_h_r_14_34257),
    .O(seg_9_5_local_g0_6_37995)
  );
  Span4Mux_h1 t3158 (
    .I(seg_8_5_sp4_v_t_38_30558),
    .O(seg_9_5_sp4_h_r_14_34257)
  );
  Span4Mux_v4 t3159 (
    .I(seg_8_9_sp4_v_t_38_31050),
    .O(seg_8_5_sp4_v_t_38_30558)
  );
  CascadeMux t316 (
    .I(net_20520),
    .O(net_20520_cascademuxed)
  );
  Span4Mux_v4 t3160 (
    .I(seg_8_13_sp4_v_t_42_31546),
    .O(seg_8_9_sp4_v_t_38_31050)
  );
  LocalMux t3161 (
    .I(seg_8_5_sp4_v_b_27_30312),
    .O(seg_8_5_local_g3_3_34185)
  );
  Span4Mux_v2 t3162 (
    .I(seg_8_7_sp4_v_t_38_30804),
    .O(seg_8_5_sp4_v_b_27_30312)
  );
  Span4Mux_v4 t3163 (
    .I(seg_8_11_sp4_v_t_42_31300),
    .O(seg_8_7_sp4_v_t_38_30804)
  );
  LocalMux t3164 (
    .I(seg_3_12_sp4_h_r_1_16590),
    .O(seg_3_12_local_g1_1_16504)
  );
  Span4Mux_h4 t3165 (
    .I(seg_7_12_sp4_v_t_36_27943),
    .O(seg_3_12_sp4_h_r_1_16590)
  );
  LocalMux t3166 (
    .I(seg_12_16_sp4_h_r_16_47105),
    .O(seg_12_16_local_g0_0_50835)
  );
  Span4Mux_h1 t3167 (
    .I(seg_11_16_sp4_h_l_40_31781),
    .O(seg_12_16_sp4_h_r_16_47105)
  );
  Span4Mux_h4 t3168 (
    .I(seg_7_16_sp4_v_b_5_27947),
    .O(seg_11_16_sp4_h_l_40_31781)
  );
  LocalMux t3169 (
    .I(seg_7_7_sp4_h_r_10_30669),
    .O(seg_7_7_local_g0_2_30575)
  );
  CascadeMux t317 (
    .I(net_20625),
    .O(net_20625_cascademuxed)
  );
  Span4Mux_h0 t3170 (
    .I(seg_7_7_sp4_v_t_40_27437),
    .O(seg_7_7_sp4_h_r_10_30669)
  );
  Span4Mux_v4 t3171 (
    .I(seg_7_11_sp4_v_t_39_27844),
    .O(seg_7_7_sp4_v_t_40_27437)
  );
  LocalMux t3172 (
    .I(seg_7_7_sp4_h_r_11_30670),
    .O(seg_7_7_local_g0_3_30576)
  );
  Span4Mux_h0 t3173 (
    .I(seg_7_7_sp4_v_t_46_27443),
    .O(seg_7_7_sp4_h_r_11_30670)
  );
  Span4Mux_v4 t3174 (
    .I(seg_7_11_sp4_v_t_45_27850),
    .O(seg_7_7_sp4_v_t_46_27443)
  );
  LocalMux t3175 (
    .I(seg_7_15_neigh_op_top_0_28093),
    .O(seg_7_15_local_g0_0_31557)
  );
  LocalMux t3176 (
    .I(seg_7_17_neigh_op_bot_2_28095),
    .O(seg_7_17_local_g0_2_31805)
  );
  LocalMux t3177 (
    .I(seg_7_17_neigh_op_bot_3_28096),
    .O(seg_7_17_local_g1_3_31814)
  );
  LocalMux t3178 (
    .I(seg_7_17_neigh_op_bot_4_28097),
    .O(seg_7_17_local_g0_4_31807)
  );
  LocalMux t3179 (
    .I(seg_7_17_neigh_op_bot_7_28100),
    .O(seg_7_17_local_g1_7_31818)
  );
  CascadeMux t318 (
    .I(net_20637),
    .O(net_20637_cascademuxed)
  );
  LocalMux t3180 (
    .I(seg_4_8_sp4_v_b_14_15865),
    .O(seg_4_8_local_g1_6_19848)
  );
  Span4Mux_v1 t3181 (
    .I(seg_4_9_sp4_v_t_37_16356),
    .O(seg_4_8_sp4_v_b_14_15865)
  );
  Span4Mux_v4 t3182 (
    .I(seg_4_13_sp4_v_t_41_16852),
    .O(seg_4_9_sp4_v_t_37_16356)
  );
  Span4Mux_v4 t3183 (
    .I(seg_4_17_sp4_h_r_11_21038),
    .O(seg_4_13_sp4_v_t_41_16852)
  );
  LocalMux t3184 (
    .I(seg_4_9_sp4_v_b_3_15865),
    .O(seg_4_9_local_g0_3_19960)
  );
  Span4Mux_v0 t3185 (
    .I(seg_4_9_sp4_v_t_37_16356),
    .O(seg_4_9_sp4_v_b_3_15865)
  );
  LocalMux t3186 (
    .I(seg_4_10_sp4_v_b_37_16356),
    .O(seg_4_10_local_g2_5_20101)
  );
  Span4Mux_v3 t3187 (
    .I(seg_4_13_sp4_v_t_41_16852),
    .O(seg_4_10_sp4_v_b_37_16356)
  );
  LocalMux t3188 (
    .I(seg_7_17_neigh_op_top_0_28297),
    .O(seg_7_17_local_g1_0_31811)
  );
  LocalMux t3189 (
    .I(seg_7_17_neigh_op_top_2_28299),
    .O(seg_7_17_local_g1_2_31813)
  );
  CascadeMux t319 (
    .I(net_20766),
    .O(net_20766_cascademuxed)
  );
  LocalMux t3190 (
    .I(seg_7_17_neigh_op_top_3_28300),
    .O(seg_7_17_local_g0_3_31806)
  );
  LocalMux t3191 (
    .I(seg_7_18_lutff_4_out_28301),
    .O(seg_7_18_local_g3_4_31954)
  );
  LocalMux t3192 (
    .I(seg_7_17_neigh_op_top_5_28302),
    .O(seg_7_17_local_g1_5_31816)
  );
  LocalMux t3193 (
    .I(seg_7_17_neigh_op_top_6_28303),
    .O(seg_7_17_local_g1_6_31817)
  );
  LocalMux t3194 (
    .I(seg_7_18_neigh_op_top_0_28399),
    .O(seg_7_18_local_g1_0_31934)
  );
  LocalMux t3195 (
    .I(seg_7_18_neigh_op_top_3_28402),
    .O(seg_7_18_local_g1_3_31937)
  );
  LocalMux t3196 (
    .I(seg_7_18_neigh_op_top_5_28404),
    .O(seg_7_18_local_g1_5_31939)
  );
  LocalMux t3197 (
    .I(seg_7_18_neigh_op_top_6_28405),
    .O(seg_7_18_local_g0_6_31932)
  );
  LocalMux t3198 (
    .I(seg_8_1_lutff_2_out_29755),
    .O(seg_8_1_local_g2_2_33644)
  );
  LocalMux t3199 (
    .I(seg_9_1_neigh_op_lft_3_29756),
    .O(seg_9_1_local_g1_3_37468)
  );
  CascadeMux t32 (
    .I(net_8131),
    .O(net_8131_cascademuxed)
  );
  CascadeMux t320 (
    .I(net_20877),
    .O(net_20877_cascademuxed)
  );
  LocalMux t3200 (
    .I(seg_9_1_neigh_op_lft_5_29758),
    .O(seg_9_1_local_g0_5_37462)
  );
  LocalMux t3201 (
    .I(seg_8_1_lutff_6_out_29759),
    .O(seg_8_1_local_g2_6_33648)
  );
  LocalMux t3202 (
    .I(seg_9_1_neigh_op_lft_7_29760),
    .O(seg_9_1_local_g0_7_37464)
  );
  LocalMux t3203 (
    .I(seg_8_2_lutff_0_out_29881),
    .O(seg_8_2_local_g3_0_33813)
  );
  LocalMux t3204 (
    .I(seg_10_2_sp4_h_r_28_33889),
    .O(seg_10_2_local_g3_4_41479)
  );
  LocalMux t3205 (
    .I(seg_13_4_sp4_h_r_5_53291),
    .O(seg_13_4_local_g0_5_53195)
  );
  Span4Mux_h0 t3206 (
    .I(seg_13_4_sp4_h_l_40_37967),
    .O(seg_13_4_sp4_h_r_5_53291)
  );
  Span4Mux_h4 t3207 (
    .I(seg_9_4_sp4_v_b_5_33771),
    .O(seg_13_4_sp4_h_l_40_37967)
  );
  LocalMux t3208 (
    .I(seg_8_3_lutff_5_out_30045),
    .O(seg_8_3_local_g0_5_33917)
  );
  LocalMux t3209 (
    .I(seg_8_3_lutff_7_out_30047),
    .O(seg_8_3_local_g2_7_33935)
  );
  CascadeMux t321 (
    .I(net_20883),
    .O(net_20883_cascademuxed)
  );
  LocalMux t3210 (
    .I(seg_7_15_sp4_v_b_10_27852),
    .O(seg_7_15_local_g1_2_31567)
  );
  Span4Mux_v4 t3211 (
    .I(seg_7_11_sp4_v_b_7_27439),
    .O(seg_7_15_sp4_v_b_10_27852)
  );
  Span4Mux_v4 t3212 (
    .I(seg_7_7_sp4_v_b_11_27035),
    .O(seg_7_11_sp4_v_b_7_27439)
  );
  Span4Mux_v4 t3213 (
    .I(seg_7_3_sp4_h_r_5_30182),
    .O(seg_7_7_sp4_v_b_11_27035)
  );
  LocalMux t3214 (
    .I(seg_8_16_sp4_v_b_21_31549),
    .O(seg_8_16_local_g1_5_35524)
  );
  Span4Mux_v3 t3215 (
    .I(seg_8_13_sp4_v_b_0_31049),
    .O(seg_8_16_sp4_v_b_21_31549)
  );
  Span4Mux_v4 t3216 (
    .I(seg_8_9_sp4_v_b_0_30557),
    .O(seg_8_13_sp4_v_b_0_31049)
  );
  Span4Mux_v4 t3217 (
    .I(seg_8_5_sp4_v_b_4_30069),
    .O(seg_8_9_sp4_v_b_0_30557)
  );
  LocalMux t3218 (
    .I(seg_8_4_lutff_2_out_30165),
    .O(seg_8_4_local_g2_2_34053)
  );
  LocalMux t3219 (
    .I(seg_7_4_neigh_op_rgt_4_30167),
    .O(seg_7_4_local_g2_4_30224)
  );
  CascadeMux t322 (
    .I(net_21006),
    .O(net_21006_cascademuxed)
  );
  LocalMux t3220 (
    .I(seg_8_4_lutff_5_out_30168),
    .O(seg_8_4_local_g0_5_34040)
  );
  LocalMux t3221 (
    .I(seg_10_3_sp4_r_v_b_16_41433),
    .O(seg_10_3_local_g3_0_41598)
  );
  Span4Mux_v1 t3222 (
    .I(seg_11_4_sp4_h_l_40_30305),
    .O(seg_10_3_sp4_r_v_b_16_41433)
  );
  LocalMux t3223 (
    .I(seg_10_3_sp4_r_v_b_22_41439),
    .O(seg_10_3_local_g3_6_41604)
  );
  Span4Mux_v1 t3224 (
    .I(seg_11_4_sp4_h_l_46_30301),
    .O(seg_10_3_sp4_r_v_b_22_41439)
  );
  LocalMux t3225 (
    .I(seg_11_1_sp4_h_r_24_37555),
    .O(seg_11_1_local_g2_0_45135)
  );
  Span4Mux_h2 t3226 (
    .I(seg_9_1_sp4_v_t_37_33896),
    .O(seg_11_1_sp4_h_r_24_37555)
  );
  LocalMux t3227 (
    .I(seg_10_3_sp4_h_r_23_37839),
    .O(seg_10_3_local_g1_7_41589)
  );
  Span4Mux_h1 t3228 (
    .I(seg_9_3_sp4_v_t_47_34152),
    .O(seg_10_3_sp4_h_r_23_37839)
  );
  LocalMux t3229 (
    .I(seg_8_5_lutff_1_out_30287),
    .O(seg_8_5_local_g1_1_34167)
  );
  CascadeMux t323 (
    .I(net_21117),
    .O(net_21117_cascademuxed)
  );
  LocalMux t3230 (
    .I(seg_7_5_neigh_op_rgt_3_30289),
    .O(seg_7_5_local_g2_3_30346)
  );
  LocalMux t3231 (
    .I(seg_8_5_lutff_4_out_30290),
    .O(seg_8_5_local_g3_4_34186)
  );
  LocalMux t3232 (
    .I(seg_8_5_lutff_5_out_30291),
    .O(seg_8_5_local_g3_5_34187)
  );
  LocalMux t3233 (
    .I(seg_7_5_neigh_op_rgt_7_30293),
    .O(seg_7_5_local_g3_7_30358)
  );
  LocalMux t3234 (
    .I(seg_8_11_sp12_v_b_0_33605),
    .O(seg_8_11_local_g3_0_34920)
  );
  LocalMux t3235 (
    .I(seg_8_9_sp4_v_b_6_30563),
    .O(seg_8_9_local_g1_6_34664)
  );
  Span4Mux_v4 t3236 (
    .I(seg_8_5_sp4_h_r_0_34252),
    .O(seg_8_9_sp4_v_b_6_30563)
  );
  LocalMux t3237 (
    .I(seg_0_7_sp4_r_v_b_34_1443),
    .O(seg_0_7_local_g2_2_1478)
  );
  Span4Mux_v2 t3238 (
    .I(seg_1_5_sp4_h_r_4_7467),
    .O(seg_0_7_sp4_r_v_b_34_1443)
  );
  Span4Mux_h4 t3239 (
    .I(seg_5_5_sp4_h_r_1_23391),
    .O(seg_1_5_sp4_h_r_4_7467)
  );
  CascadeMux t324 (
    .I(net_21222),
    .O(net_21222_cascademuxed)
  );
  LocalMux t3240 (
    .I(seg_0_17_sp4_r_v_b_1_3136),
    .O(seg_0_17_local_g1_1_3589)
  );
  Span4Mux_v4 t3241 (
    .I(seg_1_13_sp4_v_b_1_2286),
    .O(seg_0_17_sp4_r_v_b_1_3136)
  );
  Span4Mux_v4 t3242 (
    .I(seg_1_9_sp4_v_b_10_1443),
    .O(seg_1_13_sp4_v_b_1_2286)
  );
  Span4Mux_v4 t3243 (
    .I(seg_1_5_sp4_h_r_4_7467),
    .O(seg_1_9_sp4_v_b_10_1443)
  );
  LocalMux t3244 (
    .I(seg_10_19_sp4_h_r_22_39808),
    .O(seg_10_19_local_g1_6_43556)
  );
  Span4Mux_h1 t3245 (
    .I(seg_9_19_sp4_v_b_5_35621),
    .O(seg_10_19_sp4_h_r_22_39808)
  );
  Span4Mux_v4 t3246 (
    .I(seg_9_15_sp4_v_b_2_35128),
    .O(seg_9_19_sp4_v_b_5_35621)
  );
  Span4Mux_v4 t3247 (
    .I(seg_9_11_sp4_v_b_2_34636),
    .O(seg_9_15_sp4_v_b_2_35128)
  );
  Span4Mux_v4 t3248 (
    .I(seg_9_7_sp4_v_b_6_34148),
    .O(seg_9_11_sp4_v_b_2_34636)
  );
  LocalMux t3249 (
    .I(seg_7_15_sp4_r_v_b_10_31305),
    .O(seg_7_15_local_g2_2_31575)
  );
  CascadeMux t325 (
    .I(net_21258),
    .O(net_21258_cascademuxed)
  );
  Span4Mux_v4 t3250 (
    .I(seg_8_11_sp4_v_b_2_30805),
    .O(seg_7_15_sp4_r_v_b_10_31305)
  );
  Span4Mux_v4 t3251 (
    .I(seg_8_7_sp4_v_b_11_30320),
    .O(seg_8_11_sp4_v_b_2_30805)
  );
  LocalMux t3252 (
    .I(seg_7_15_sp4_r_v_b_21_31426),
    .O(seg_7_15_local_g3_5_31586)
  );
  Span4Mux_v3 t3253 (
    .I(seg_8_12_sp4_v_b_5_30929),
    .O(seg_7_15_sp4_r_v_b_21_31426)
  );
  Span4Mux_v4 t3254 (
    .I(seg_8_8_sp4_v_b_2_30436),
    .O(seg_8_12_sp4_v_b_5_30929)
  );
  LocalMux t3255 (
    .I(seg_7_15_sp4_r_v_b_20_31425),
    .O(seg_7_15_local_g3_4_31585)
  );
  Span4Mux_v3 t3256 (
    .I(seg_8_12_sp4_v_b_9_30933),
    .O(seg_7_15_sp4_r_v_b_20_31425)
  );
  Span4Mux_v4 t3257 (
    .I(seg_8_8_sp4_v_b_6_30440),
    .O(seg_8_12_sp4_v_b_9_30933)
  );
  LocalMux t3258 (
    .I(seg_7_15_sp4_r_v_b_17_31422),
    .O(seg_7_15_local_g3_1_31582)
  );
  Span4Mux_v3 t3259 (
    .I(seg_8_12_sp4_v_b_4_30930),
    .O(seg_7_15_sp4_r_v_b_17_31422)
  );
  CascadeMux t326 (
    .I(net_21264),
    .O(net_21264_cascademuxed)
  );
  Span4Mux_v4 t3260 (
    .I(seg_8_8_sp4_v_b_8_30442),
    .O(seg_8_12_sp4_v_b_4_30930)
  );
  LocalMux t3261 (
    .I(seg_8_16_sp4_v_b_16_31544),
    .O(seg_8_16_local_g1_0_35519)
  );
  Span4Mux_v3 t3262 (
    .I(seg_8_13_sp4_v_b_5_31052),
    .O(seg_8_16_sp4_v_b_16_31544)
  );
  Span4Mux_v4 t3263 (
    .I(seg_8_9_sp4_v_b_5_30560),
    .O(seg_8_13_sp4_v_b_5_31052)
  );
  LocalMux t3264 (
    .I(seg_8_16_sp4_v_b_20_31548),
    .O(seg_8_16_local_g0_4_35515)
  );
  Span4Mux_v3 t3265 (
    .I(seg_8_13_sp4_v_b_9_31056),
    .O(seg_8_16_sp4_v_b_20_31548)
  );
  Span4Mux_v4 t3266 (
    .I(seg_8_9_sp4_v_b_9_30564),
    .O(seg_8_13_sp4_v_b_9_31056)
  );
  LocalMux t3267 (
    .I(seg_8_16_sp12_v_b_3_34251),
    .O(seg_8_16_local_g2_3_35530)
  );
  LocalMux t3268 (
    .I(seg_8_16_sp4_r_v_b_16_35375),
    .O(seg_8_16_local_g3_0_35535)
  );
  Span4Mux_v3 t3269 (
    .I(seg_9_13_sp4_v_b_5_34883),
    .O(seg_8_16_sp4_r_v_b_16_35375)
  );
  CascadeMux t327 (
    .I(net_21375),
    .O(net_21375_cascademuxed)
  );
  Span4Mux_v4 t3270 (
    .I(seg_9_9_sp4_v_b_5_34391),
    .O(seg_9_13_sp4_v_b_5_34883)
  );
  LocalMux t3271 (
    .I(seg_8_16_sp4_v_b_15_31543),
    .O(seg_8_16_local_g1_7_35526)
  );
  Span4Mux_v3 t3272 (
    .I(seg_8_13_sp4_v_b_11_31058),
    .O(seg_8_16_sp4_v_b_15_31543)
  );
  Span4Mux_v4 t3273 (
    .I(seg_8_9_sp4_v_b_8_30565),
    .O(seg_8_13_sp4_v_b_11_31058)
  );
  LocalMux t3274 (
    .I(seg_9_8_neigh_op_lft_1_30656),
    .O(seg_9_8_local_g0_1_38359)
  );
  LocalMux t3275 (
    .I(seg_9_8_neigh_op_lft_2_30657),
    .O(seg_9_8_local_g1_2_38368)
  );
  LocalMux t3276 (
    .I(seg_9_8_neigh_op_lft_3_30658),
    .O(seg_9_8_local_g0_3_38361)
  );
  LocalMux t3277 (
    .I(seg_9_8_neigh_op_lft_4_30659),
    .O(seg_9_8_local_g1_4_38370)
  );
  LocalMux t3278 (
    .I(seg_9_8_neigh_op_lft_5_30660),
    .O(seg_9_8_local_g0_5_38363)
  );
  LocalMux t3279 (
    .I(seg_9_8_neigh_op_lft_6_30661),
    .O(seg_9_8_local_g0_6_38364)
  );
  CascadeMux t328 (
    .I(net_22817),
    .O(net_22817_cascademuxed)
  );
  LocalMux t3280 (
    .I(seg_9_8_neigh_op_lft_7_30662),
    .O(seg_9_8_local_g0_7_38365)
  );
  LocalMux t3281 (
    .I(seg_9_8_neigh_op_tnl_1_30779),
    .O(seg_9_8_local_g2_1_38375)
  );
  LocalMux t3282 (
    .I(seg_8_9_lutff_2_out_30780),
    .O(seg_8_9_local_g0_2_34652)
  );
  LocalMux t3283 (
    .I(seg_8_8_neigh_op_top_4_30782),
    .O(seg_8_8_local_g1_4_34539)
  );
  LocalMux t3284 (
    .I(seg_8_9_lutff_4_out_30782),
    .O(seg_8_9_local_g1_4_34662)
  );
  LocalMux t3285 (
    .I(seg_8_8_neigh_op_top_5_30783),
    .O(seg_8_8_local_g1_5_34540)
  );
  LocalMux t3286 (
    .I(seg_8_9_lutff_6_out_30784),
    .O(seg_8_9_local_g2_6_34672)
  );
  LocalMux t3287 (
    .I(seg_8_8_neigh_op_top_7_30785),
    .O(seg_8_8_local_g1_7_34542)
  );
  LocalMux t3288 (
    .I(seg_8_9_lutff_7_out_30785),
    .O(seg_8_9_local_g1_7_34665)
  );
  LocalMux t3289 (
    .I(seg_8_4_sp4_r_v_b_12_33895),
    .O(seg_8_4_local_g2_4_34055)
  );
  CascadeMux t329 (
    .I(net_22841),
    .O(net_22841_cascademuxed)
  );
  Span4Mux_v1 t3290 (
    .I(seg_9_5_sp4_v_t_36_34387),
    .O(seg_8_4_sp4_r_v_b_12_33895)
  );
  LocalMux t3291 (
    .I(seg_8_15_sp4_v_b_12_31417),
    .O(seg_8_15_local_g0_4_35392)
  );
  Span4Mux_v3 t3292 (
    .I(seg_8_12_sp4_v_b_10_30936),
    .O(seg_8_15_sp4_v_b_12_31417)
  );
  LocalMux t3293 (
    .I(seg_8_15_sp4_v_b_25_31540),
    .O(seg_8_15_local_g3_1_35413)
  );
  Span4Mux_v2 t3294 (
    .I(seg_8_13_sp4_v_b_1_31048),
    .O(seg_8_15_sp4_v_b_25_31540)
  );
  LocalMux t3295 (
    .I(seg_8_11_lutff_0_out_31024),
    .O(seg_8_11_local_g1_0_34904)
  );
  LocalMux t3296 (
    .I(seg_7_12_neigh_op_bnr_1_31025),
    .O(seg_7_12_local_g1_1_31197)
  );
  LocalMux t3297 (
    .I(seg_8_11_lutff_2_out_31026),
    .O(seg_8_11_local_g1_2_34906)
  );
  LocalMux t3298 (
    .I(seg_7_12_neigh_op_bnr_3_31027),
    .O(seg_7_12_local_g0_3_31191)
  );
  LocalMux t3299 (
    .I(seg_9_12_neigh_op_bnl_3_31027),
    .O(seg_9_12_local_g3_3_38877)
  );
  CascadeMux t33 (
    .I(net_8143),
    .O(net_8143_cascademuxed)
  );
  CascadeMux t330 (
    .I(net_22968),
    .O(net_22968_cascademuxed)
  );
  LocalMux t3300 (
    .I(seg_9_10_neigh_op_tnl_4_31028),
    .O(seg_9_10_local_g3_4_38632)
  );
  LocalMux t3301 (
    .I(seg_8_11_lutff_6_out_31030),
    .O(seg_8_11_local_g2_6_34918)
  );
  LocalMux t3302 (
    .I(seg_14_10_sp4_r_v_b_16_57622),
    .O(seg_14_10_local_g3_0_57782)
  );
  Span4Mux_v1 t3303 (
    .I(seg_15_11_sp4_h_l_46_46486),
    .O(seg_14_10_sp4_r_v_b_16_57622)
  );
  Span4Mux_h4 t3304 (
    .I(seg_11_11_sp4_h_l_38_31164),
    .O(seg_15_11_sp4_h_l_46_46486)
  );
  LocalMux t3305 (
    .I(seg_8_6_sp4_r_v_b_29_34268),
    .O(seg_8_6_local_g1_5_34294)
  );
  Span4Mux_v2 t3306 (
    .I(seg_9_8_sp4_v_t_39_34759),
    .O(seg_8_6_sp4_r_v_b_29_34268)
  );
  LocalMux t3307 (
    .I(seg_9_4_sp4_h_r_10_37962),
    .O(seg_9_4_local_g1_2_37876)
  );
  Span4Mux_h0 t3308 (
    .I(seg_9_4_sp4_v_t_40_34268),
    .O(seg_9_4_sp4_h_r_10_37962)
  );
  Span4Mux_v4 t3309 (
    .I(seg_9_8_sp4_v_t_39_34759),
    .O(seg_9_4_sp4_v_t_40_34268)
  );
  CascadeMux t331 (
    .I(net_23127),
    .O(net_23127_cascademuxed)
  );
  LocalMux t3310 (
    .I(seg_10_4_sp4_h_r_23_37962),
    .O(seg_10_4_local_g0_7_41704)
  );
  Span4Mux_h1 t3311 (
    .I(seg_9_4_sp4_v_t_40_34268),
    .O(seg_10_4_sp4_h_r_23_37962)
  );
  LocalMux t3312 (
    .I(seg_8_8_sp4_v_b_47_30813),
    .O(seg_8_8_local_g3_7_34558)
  );
  LocalMux t3313 (
    .I(seg_7_9_sp4_r_v_b_38_30927),
    .O(seg_7_9_local_g2_6_30841)
  );
  LocalMux t3314 (
    .I(seg_9_8_sp4_v_b_23_34398),
    .O(seg_9_8_local_g1_7_38373)
  );
  Span4Mux_v1 t3315 (
    .I(seg_9_9_sp4_v_t_39_34882),
    .O(seg_9_8_sp4_v_b_23_34398)
  );
  LocalMux t3316 (
    .I(seg_8_13_lutff_0_out_31270),
    .O(seg_8_13_local_g2_0_35158)
  );
  LocalMux t3317 (
    .I(seg_7_12_neigh_op_tnr_3_31273),
    .O(seg_7_12_local_g2_3_31207)
  );
  LocalMux t3318 (
    .I(seg_8_13_lutff_4_out_31274),
    .O(seg_8_13_local_g1_4_35154)
  );
  LocalMux t3319 (
    .I(seg_7_12_neigh_op_tnr_5_31275),
    .O(seg_7_12_local_g3_5_31217)
  );
  CascadeMux t332 (
    .I(net_23220),
    .O(net_23220_cascademuxed)
  );
  LocalMux t3320 (
    .I(seg_9_12_neigh_op_tnl_5_31275),
    .O(seg_9_12_local_g3_5_38879)
  );
  LocalMux t3321 (
    .I(seg_8_13_lutff_6_out_31276),
    .O(seg_8_13_local_g3_6_35172)
  );
  LocalMux t3322 (
    .I(seg_9_8_sp4_v_b_38_34635),
    .O(seg_9_8_local_g2_6_38380)
  );
  Span4Mux_v3 t3323 (
    .I(seg_9_11_sp4_v_t_42_35131),
    .O(seg_9_8_sp4_v_b_38_34635)
  );
  LocalMux t3324 (
    .I(seg_8_11_sp4_v_b_26_31051),
    .O(seg_8_11_local_g3_2_34922)
  );
  LocalMux t3325 (
    .I(seg_8_4_sp4_v_b_18_30070),
    .O(seg_8_4_local_g1_2_34045)
  );
  Span4Mux_v1 t3326 (
    .I(seg_8_5_sp4_v_t_41_30561),
    .O(seg_8_4_sp4_v_b_18_30070)
  );
  Span4Mux_v4 t3327 (
    .I(seg_8_9_sp4_v_t_41_31053),
    .O(seg_8_5_sp4_v_t_41_30561)
  );
  LocalMux t3328 (
    .I(seg_8_14_lutff_0_out_31393),
    .O(seg_8_14_local_g2_0_35281)
  );
  LocalMux t3329 (
    .I(seg_7_15_neigh_op_bnr_6_31399),
    .O(seg_7_15_local_g1_6_31571)
  );
  CascadeMux t333 (
    .I(net_23232),
    .O(net_23232_cascademuxed)
  );
  LocalMux t3330 (
    .I(seg_12_14_sp4_v_b_19_46625),
    .O(seg_12_14_local_g1_3_50600)
  );
  Span4Mux_v1 t3331 (
    .I(seg_12_15_sp4_h_l_37_35482),
    .O(seg_12_14_sp4_v_b_19_46625)
  );
  LocalMux t3332 (
    .I(seg_10_18_sp4_r_v_b_12_43279),
    .O(seg_10_18_local_g2_4_43439)
  );
  Span4Mux_v3 t3333 (
    .I(seg_11_15_sp4_h_l_36_31652),
    .O(seg_10_18_sp4_r_v_b_12_43279)
  );
  LocalMux t3334 (
    .I(seg_12_14_sp4_v_b_17_46623),
    .O(seg_12_14_local_g0_1_50590)
  );
  Span4Mux_v1 t3335 (
    .I(seg_12_15_sp4_h_l_41_35488),
    .O(seg_12_14_sp4_v_b_17_46623)
  );
  LocalMux t3336 (
    .I(seg_11_12_sp4_h_r_31_38953),
    .O(seg_11_12_local_g2_7_46535)
  );
  Span4Mux_h2 t3337 (
    .I(seg_9_12_sp4_v_t_39_35251),
    .O(seg_11_12_sp4_h_r_31_38953)
  );
  LocalMux t3338 (
    .I(seg_13_8_sp4_v_b_44_49965),
    .O(seg_13_8_local_g2_4_53702)
  );
  Span4Mux_v3 t3339 (
    .I(seg_13_11_sp4_h_l_38_38826),
    .O(seg_13_8_sp4_v_b_44_49965)
  );
  CascadeMux t334 (
    .I(net_23331),
    .O(net_23331_cascademuxed)
  );
  Span4Mux_h4 t3340 (
    .I(seg_9_11_sp4_v_t_38_35127),
    .O(seg_13_11_sp4_h_l_38_38826)
  );
  LocalMux t3341 (
    .I(seg_12_14_sp4_h_r_39_39194),
    .O(seg_12_14_local_g2_7_50612)
  );
  Span4Mux_h3 t3342 (
    .I(seg_9_14_sp4_v_t_39_35497),
    .O(seg_12_14_sp4_h_r_39_39194)
  );
  LocalMux t3343 (
    .I(seg_12_14_sp4_h_r_44_39201),
    .O(seg_12_14_local_g2_4_50609)
  );
  Span4Mux_h3 t3344 (
    .I(seg_9_14_sp4_v_t_41_35499),
    .O(seg_12_14_sp4_h_r_44_39201)
  );
  LocalMux t3345 (
    .I(seg_9_5_sp4_h_r_0_38083),
    .O(seg_9_5_local_g1_0_37997)
  );
  Span4Mux_h0 t3346 (
    .I(seg_9_5_sp4_v_t_37_34388),
    .O(seg_9_5_sp4_h_r_0_38083)
  );
  Span4Mux_v4 t3347 (
    .I(seg_9_9_sp4_v_t_37_34880),
    .O(seg_9_5_sp4_v_t_37_34388)
  );
  Span4Mux_v4 t3348 (
    .I(seg_9_13_sp4_v_t_37_35372),
    .O(seg_9_9_sp4_v_t_37_34880)
  );
  LocalMux t3349 (
    .I(seg_9_10_sp4_v_b_44_34887),
    .O(seg_9_10_local_g2_4_38624)
  );
  CascadeMux t335 (
    .I(net_23361),
    .O(net_23361_cascademuxed)
  );
  Span4Mux_v3 t3350 (
    .I(seg_9_13_sp4_v_t_43_35378),
    .O(seg_9_10_sp4_v_b_44_34887)
  );
  LocalMux t3351 (
    .I(seg_8_9_sp4_r_v_b_42_34762),
    .O(seg_8_9_local_g3_2_34676)
  );
  Span4Mux_v3 t3352 (
    .I(seg_9_12_sp4_v_t_42_35254),
    .O(seg_8_9_sp4_r_v_b_42_34762)
  );
  LocalMux t3353 (
    .I(seg_3_3_sp4_r_v_b_28_15376),
    .O(seg_3_3_local_g1_4_15400)
  );
  Span4Mux_v2 t3354 (
    .I(seg_4_5_sp4_h_r_4_19565),
    .O(seg_3_3_sp4_r_v_b_28_15376)
  );
  Span4Mux_h4 t3355 (
    .I(seg_8_5_sp4_v_t_47_30567),
    .O(seg_4_5_sp4_h_r_4_19565)
  );
  Sp12to4 t3356 (
    .I(seg_8_8_sp12_v_b_23_34497),
    .O(seg_8_5_sp4_v_t_47_30567)
  );
  Span12Mux_v11 t3357 (
    .I(seg_8_19_sp12_v_t_23_35973),
    .O(seg_8_8_sp12_v_b_23_34497)
  );
  LocalMux t3358 (
    .I(seg_4_3_sp4_v_b_28_15376),
    .O(seg_4_3_local_g2_4_19239)
  );
  Span4Mux_v2 t3359 (
    .I(seg_4_5_sp4_h_r_4_19565),
    .O(seg_4_3_sp4_v_b_28_15376)
  );
  CascadeMux t336 (
    .I(net_23454),
    .O(net_23454_cascademuxed)
  );
  LocalMux t3360 (
    .I(seg_3_2_sp4_r_v_b_44_15379),
    .O(seg_3_2_local_g3_4_15293)
  );
  Span4Mux_v3 t3361 (
    .I(seg_4_5_sp4_v_t_36_15863),
    .O(seg_3_2_sp4_r_v_b_44_15379)
  );
  Span4Mux_v4 t3362 (
    .I(seg_4_9_sp4_h_r_8_20061),
    .O(seg_4_5_sp4_v_t_36_15863)
  );
  Span4Mux_h4 t3363 (
    .I(seg_8_9_sp4_v_t_45_31057),
    .O(seg_4_9_sp4_h_r_8_20061)
  );
  Sp12to4 t3364 (
    .I(seg_8_12_sp12_v_b_19_34743),
    .O(seg_8_9_sp4_v_t_45_31057)
  );
  Span12Mux_v9 t3365 (
    .I(seg_8_21_sp12_v_t_23_36219),
    .O(seg_8_12_sp12_v_b_19_34743)
  );
  LocalMux t3366 (
    .I(seg_4_2_sp4_v_b_44_15379),
    .O(seg_4_2_local_g3_4_19124)
  );
  Span4Mux_v3 t3367 (
    .I(seg_4_5_sp4_v_t_36_15863),
    .O(seg_4_2_sp4_v_b_44_15379)
  );
  LocalMux t3368 (
    .I(seg_10_1_neigh_op_lft_1_33585),
    .O(seg_10_1_local_g0_1_41289)
  );
  LocalMux t3369 (
    .I(seg_10_1_neigh_op_lft_3_33587),
    .O(seg_10_1_local_g1_3_41299)
  );
  CascadeMux t337 (
    .I(net_23460),
    .O(net_23460_cascademuxed)
  );
  LocalMux t3370 (
    .I(seg_10_1_neigh_op_lft_4_33588),
    .O(seg_10_1_local_g0_4_41292)
  );
  LocalMux t3371 (
    .I(seg_10_1_neigh_op_lft_6_33590),
    .O(seg_10_1_local_g1_6_41302)
  );
  LocalMux t3372 (
    .I(seg_9_1_lutff_7_out_33591),
    .O(seg_9_1_local_g2_7_37480)
  );
  LocalMux t3373 (
    .I(seg_9_3_neigh_op_bot_3_33715),
    .O(seg_9_3_local_g0_3_37746)
  );
  LocalMux t3374 (
    .I(seg_8_3_neigh_op_bnr_6_33718),
    .O(seg_8_3_local_g0_6_33918)
  );
  LocalMux t3375 (
    .I(seg_9_3_lutff_3_out_33874),
    .O(seg_9_3_local_g2_3_37762)
  );
  LocalMux t3376 (
    .I(seg_8_16_sp4_r_v_b_14_35373),
    .O(seg_8_16_local_g2_6_35533)
  );
  Span4Mux_v3 t3377 (
    .I(seg_9_13_sp4_v_b_7_34885),
    .O(seg_8_16_sp4_r_v_b_14_35373)
  );
  Span4Mux_v4 t3378 (
    .I(seg_9_9_sp4_v_b_4_34392),
    .O(seg_9_13_sp4_v_b_7_34885)
  );
  Span4Mux_v4 t3379 (
    .I(seg_9_5_sp4_v_b_4_33900),
    .O(seg_9_9_sp4_v_b_4_34392)
  );
  CascadeMux t338 (
    .I(net_23466),
    .O(net_23466_cascademuxed)
  );
  LocalMux t3380 (
    .I(seg_9_4_lutff_2_out_33996),
    .O(seg_9_4_local_g2_2_37884)
  );
  LocalMux t3381 (
    .I(seg_10_4_neigh_op_lft_6_34000),
    .O(seg_10_4_local_g0_6_41703)
  );
  LocalMux t3382 (
    .I(seg_10_4_neigh_op_lft_7_34001),
    .O(seg_10_4_local_g1_7_41712)
  );
  LocalMux t3383 (
    .I(seg_7_5_sp4_v_b_45_27136),
    .O(seg_7_5_local_g2_5_30348)
  );
  Span4Mux_v1 t3384 (
    .I(seg_7_4_sp4_h_r_2_30302),
    .O(seg_7_5_sp4_v_b_45_27136)
  );
  LocalMux t3385 (
    .I(seg_7_15_sp4_v_b_23_27954),
    .O(seg_7_15_local_g0_7_31564)
  );
  Span4Mux_v3 t3386 (
    .I(seg_7_12_sp4_v_b_10_27546),
    .O(seg_7_15_sp4_v_b_23_27954)
  );
  Span4Mux_v4 t3387 (
    .I(seg_7_8_sp4_v_b_2_27130),
    .O(seg_7_12_sp4_v_b_10_27546)
  );
  Span4Mux_v4 t3388 (
    .I(seg_7_4_sp4_h_r_8_30308),
    .O(seg_7_8_sp4_v_b_2_27130)
  );
  LocalMux t3389 (
    .I(seg_10_5_neigh_op_lft_0_34117),
    .O(seg_10_5_local_g1_0_41828)
  );
  CascadeMux t339 (
    .I(net_23472),
    .O(net_23472_cascademuxed)
  );
  LocalMux t3390 (
    .I(seg_9_5_lutff_3_out_34120),
    .O(seg_9_5_local_g3_3_38016)
  );
  LocalMux t3391 (
    .I(seg_9_5_lutff_6_out_34123),
    .O(seg_9_5_local_g2_6_38011)
  );
  LocalMux t3392 (
    .I(seg_7_5_sp4_h_r_10_30423),
    .O(seg_7_5_local_g0_2_30329)
  );
  LocalMux t3393 (
    .I(seg_7_5_sp4_h_r_22_27118),
    .O(seg_7_5_local_g0_6_30333)
  );
  LocalMux t3394 (
    .I(seg_9_1_sp4_h_r_8_37565),
    .O(seg_9_1_local_g0_0_37457)
  );
  Span4Mux_h0 t3395 (
    .I(seg_9_1_sp4_v_t_45_33904),
    .O(seg_9_1_sp4_h_r_8_37565)
  );
  LocalMux t3396 (
    .I(seg_9_6_lutff_0_out_34240),
    .O(seg_9_6_local_g1_0_38120)
  );
  LocalMux t3397 (
    .I(seg_10_5_neigh_op_tnl_2_34242),
    .O(seg_10_5_local_g3_2_41846)
  );
  LocalMux t3398 (
    .I(seg_11_6_sp4_h_r_46_34378),
    .O(seg_11_6_local_g2_6_45796)
  );
  LocalMux t3399 (
    .I(seg_10_2_sp4_h_r_9_41556),
    .O(seg_10_2_local_g0_1_41452)
  );
  CascadeMux t34 (
    .I(net_8149),
    .O(net_8149_cascademuxed)
  );
  CascadeMux t340 (
    .I(net_23478),
    .O(net_23478_cascademuxed)
  );
  Span4Mux_h0 t3400 (
    .I(seg_10_2_sp4_v_t_44_37857),
    .O(seg_10_2_sp4_h_r_9_41556)
  );
  LocalMux t3401 (
    .I(seg_10_7_neigh_op_lft_0_34363),
    .O(seg_10_7_local_g1_0_42074)
  );
  LocalMux t3402 (
    .I(seg_8_6_neigh_op_tnr_1_34364),
    .O(seg_8_6_local_g2_1_34298)
  );
  LocalMux t3403 (
    .I(seg_9_7_lutff_2_out_34365),
    .O(seg_9_7_local_g2_2_38253)
  );
  LocalMux t3404 (
    .I(seg_9_7_lutff_3_out_34366),
    .O(seg_9_7_local_g1_3_38246)
  );
  LocalMux t3405 (
    .I(seg_9_7_lutff_4_out_34367),
    .O(seg_9_7_local_g2_4_38255)
  );
  LocalMux t3406 (
    .I(seg_9_7_lutff_6_out_34369),
    .O(seg_9_7_local_g1_6_38249)
  );
  LocalMux t3407 (
    .I(seg_9_6_neigh_op_top_7_34370),
    .O(seg_9_6_local_g1_7_38127)
  );
  LocalMux t3408 (
    .I(seg_0_25_sp12_v_b_13_4134),
    .O(seg_0_25_local_g2_5_5342)
  );
  Span12Mux_v6 t3409 (
    .I(seg_0_19_sp12_v_b_1_1578),
    .O(seg_0_25_sp12_v_b_13_4134)
  );
  CascadeMux t341 (
    .I(net_23484),
    .O(net_23484_cascademuxed)
  );
  Span12Mux_v12 t3410 (
    .I(seg_0_7_sp12_h_r_1_1555),
    .O(seg_0_19_sp12_v_b_1_1578)
  );
  LocalMux t3411 (
    .I(seg_0_12_sp12_h_r_6_2634),
    .O(seg_0_12_local_g1_6_2534)
  );
  Span12Mux_h9 t3412 (
    .I(seg_9_12_sp12_v_b_1_37438),
    .O(seg_0_12_sp12_h_r_6_2634)
  );
  LocalMux t3413 (
    .I(seg_8_14_sp4_v_b_12_31294),
    .O(seg_8_14_local_g0_4_35269)
  );
  Span4Mux_v3 t3414 (
    .I(seg_8_11_sp4_v_b_1_30802),
    .O(seg_8_14_sp4_v_b_12_31294)
  );
  Span4Mux_v4 t3415 (
    .I(seg_8_7_sp4_h_r_7_34507),
    .O(seg_8_11_sp4_v_b_1_30802)
  );
  LocalMux t3416 (
    .I(seg_14_6_sp4_v_b_20_53304),
    .O(seg_14_6_local_g1_4_57278)
  );
  Span4Mux_v1 t3417 (
    .I(seg_14_7_sp4_h_l_38_42165),
    .O(seg_14_6_sp4_v_b_20_53304)
  );
  Span4Mux_h4 t3418 (
    .I(seg_10_7_sp4_v_b_3_37974),
    .O(seg_14_7_sp4_h_l_38_42165)
  );
  LocalMux t3419 (
    .I(seg_7_9_sp4_h_r_17_27529),
    .O(seg_7_9_local_g0_1_30820)
  );
  CascadeMux t342 (
    .I(net_23496),
    .O(net_23496_cascademuxed)
  );
  Span4Mux_h3 t3420 (
    .I(seg_10_9_sp4_v_b_11_38228),
    .O(seg_7_9_sp4_h_r_17_27529)
  );
  LocalMux t3421 (
    .I(seg_10_12_sp4_v_b_18_38716),
    .O(seg_10_12_local_g0_2_42683)
  );
  Span4Mux_v3 t3422 (
    .I(seg_10_9_sp4_v_b_11_38228),
    .O(seg_10_12_sp4_v_b_18_38716)
  );
  LocalMux t3423 (
    .I(seg_9_7_neigh_op_top_1_34487),
    .O(seg_9_7_local_g1_1_38244)
  );
  LocalMux t3424 (
    .I(seg_10_8_neigh_op_lft_2_34488),
    .O(seg_10_8_local_g1_2_42199)
  );
  LocalMux t3425 (
    .I(seg_10_7_neigh_op_tnl_3_34489),
    .O(seg_10_7_local_g3_3_42093)
  );
  LocalMux t3426 (
    .I(seg_10_8_neigh_op_lft_4_34490),
    .O(seg_10_8_local_g0_4_42193)
  );
  LocalMux t3427 (
    .I(seg_10_8_neigh_op_lft_5_34491),
    .O(seg_10_8_local_g1_5_42202)
  );
  LocalMux t3428 (
    .I(seg_10_8_neigh_op_lft_6_34492),
    .O(seg_10_8_local_g1_6_42203)
  );
  LocalMux t3429 (
    .I(seg_11_4_sp4_h_r_5_45629),
    .O(seg_11_4_local_g0_5_45533)
  );
  CascadeMux t343 (
    .I(net_23583),
    .O(net_23583_cascademuxed)
  );
  Span4Mux_h0 t3430 (
    .I(seg_11_4_sp4_v_t_37_41927),
    .O(seg_11_4_sp4_h_r_5_45629)
  );
  Span4Mux_v4 t3431 (
    .I(seg_11_8_sp4_h_l_43_30798),
    .O(seg_11_4_sp4_v_t_37_41927)
  );
  LocalMux t3432 (
    .I(seg_13_3_sp4_v_b_33_49227),
    .O(seg_13_3_local_g3_1_53092)
  );
  Span4Mux_v2 t3433 (
    .I(seg_13_5_sp4_h_l_38_38088),
    .O(seg_13_3_sp4_v_b_33_49227)
  );
  Span4Mux_h4 t3434 (
    .I(seg_9_5_sp4_v_t_38_34389),
    .O(seg_13_5_sp4_h_l_38_38088)
  );
  LocalMux t3435 (
    .I(seg_10_8_neigh_op_tnl_0_34609),
    .O(seg_10_8_local_g3_0_42213)
  );
  LocalMux t3436 (
    .I(seg_8_8_neigh_op_tnr_1_34610),
    .O(seg_8_8_local_g3_1_34552)
  );
  LocalMux t3437 (
    .I(seg_8_8_neigh_op_tnr_2_34611),
    .O(seg_8_8_local_g3_2_34553)
  );
  LocalMux t3438 (
    .I(seg_9_9_lutff_3_out_34612),
    .O(seg_9_9_local_g0_3_38484)
  );
  LocalMux t3439 (
    .I(seg_8_8_neigh_op_tnr_4_34613),
    .O(seg_8_8_local_g2_4_34547)
  );
  CascadeMux t344 (
    .I(net_23589),
    .O(net_23589_cascademuxed)
  );
  LocalMux t3440 (
    .I(seg_9_9_lutff_5_out_34614),
    .O(seg_9_9_local_g1_5_38494)
  );
  LocalMux t3441 (
    .I(seg_9_6_sp4_h_r_6_38214),
    .O(seg_9_6_local_g0_6_38118)
  );
  Span4Mux_h0 t3442 (
    .I(seg_9_6_sp4_v_t_36_34510),
    .O(seg_9_6_sp4_h_r_6_38214)
  );
  LocalMux t3443 (
    .I(seg_9_6_sp4_v_b_15_34144),
    .O(seg_9_6_local_g0_7_38119)
  );
  Span4Mux_v1 t3444 (
    .I(seg_9_7_sp4_v_t_43_34640),
    .O(seg_9_6_sp4_v_b_15_34144)
  );
  LocalMux t3445 (
    .I(seg_9_10_lutff_1_out_34733),
    .O(seg_9_10_local_g3_1_38629)
  );
  LocalMux t3446 (
    .I(seg_9_9_neigh_op_top_2_34734),
    .O(seg_9_9_local_g1_2_38491)
  );
  LocalMux t3447 (
    .I(seg_9_10_lutff_4_out_34736),
    .O(seg_9_10_local_g0_4_38608)
  );
  LocalMux t3448 (
    .I(seg_9_9_neigh_op_top_5_34737),
    .O(seg_9_9_local_g0_5_38486)
  );
  LocalMux t3449 (
    .I(seg_9_9_neigh_op_top_6_34738),
    .O(seg_9_9_local_g1_6_38495)
  );
  CascadeMux t345 (
    .I(net_23595),
    .O(net_23595_cascademuxed)
  );
  LocalMux t3450 (
    .I(seg_0_12_sp4_h_r_28_2673),
    .O(seg_0_12_local_g3_4_2548)
  );
  Span4Mux_h2 t3451 (
    .I(seg_2_12_sp4_h_r_8_12768),
    .O(seg_0_12_sp4_h_r_28_2673)
  );
  Span4Mux_h4 t3452 (
    .I(seg_6_12_sp4_h_r_0_27829),
    .O(seg_2_12_sp4_h_r_8_12768)
  );
  Span4Mux_h4 t3453 (
    .I(seg_10_12_sp4_v_b_7_38593),
    .O(seg_6_12_sp4_h_r_0_27829)
  );
  LocalMux t3454 (
    .I(seg_9_7_sp4_v_b_37_34511),
    .O(seg_9_7_local_g2_5_38256)
  );
  LocalMux t3455 (
    .I(seg_0_25_sp4_r_v_b_0_4878),
    .O(seg_0_25_local_g1_0_5329)
  );
  Span4Mux_v4 t3456 (
    .I(seg_1_21_sp4_v_b_0_3970),
    .O(seg_0_25_sp4_r_v_b_0_4878)
  );
  Span4Mux_v4 t3457 (
    .I(seg_1_17_sp4_h_r_0_9225),
    .O(seg_1_21_sp4_v_b_0_3970)
  );
  Span4Mux_h4 t3458 (
    .I(seg_5_17_sp4_h_r_0_24866),
    .O(seg_1_17_sp4_h_r_0_9225)
  );
  Span4Mux_h4 t3459 (
    .I(seg_9_17_sp4_v_b_7_35377),
    .O(seg_5_17_sp4_h_r_0_24866)
  );
  CascadeMux t346 (
    .I(net_23607),
    .O(net_23607_cascademuxed)
  );
  Span4Mux_v4 t3460 (
    .I(seg_9_13_sp4_v_b_11_34889),
    .O(seg_9_17_sp4_v_b_7_35377)
  );
  LocalMux t3461 (
    .I(seg_9_11_lutff_0_out_34855),
    .O(seg_9_11_local_g1_0_38735)
  );
  LocalMux t3462 (
    .I(seg_9_11_lutff_6_out_34861),
    .O(seg_9_11_local_g2_6_38749)
  );
  LocalMux t3463 (
    .I(seg_3_18_sp4_r_v_b_18_17099),
    .O(seg_3_18_local_g3_2_17259)
  );
  Span4Mux_v3 t3464 (
    .I(seg_4_15_sp4_v_b_4_16606),
    .O(seg_3_18_sp4_r_v_b_18_17099)
  );
  Span4Mux_v4 t3465 (
    .I(seg_4_11_sp4_h_r_4_20303),
    .O(seg_4_15_sp4_v_b_4_16606)
  );
  Span4Mux_h4 t3466 (
    .I(seg_8_11_sp4_h_r_1_34991),
    .O(seg_4_11_sp4_h_r_4_20303)
  );
  LocalMux t3467 (
    .I(seg_15_6_sp4_r_v_b_18_60962),
    .O(seg_15_6_local_g3_2_61122)
  );
  Span4Mux_v1 t3468 (
    .I(seg_16_7_sp4_h_l_36_49823),
    .O(seg_15_6_sp4_r_v_b_18_60962)
  );
  Span4Mux_h4 t3469 (
    .I(seg_12_7_sp4_v_t_36_46126),
    .O(seg_16_7_sp4_h_l_36_49823)
  );
  CascadeMux t347 (
    .I(net_23700),
    .O(net_23700_cascademuxed)
  );
  Span4Mux_v4 t3470 (
    .I(seg_12_11_sp4_h_l_36_34991),
    .O(seg_12_7_sp4_v_t_36_46126)
  );
  LocalMux t3471 (
    .I(seg_15_18_sp4_r_v_b_17_62437),
    .O(seg_15_18_local_g3_1_62597)
  );
  Span4Mux_v3 t3472 (
    .I(seg_16_15_sp4_v_b_1_61940),
    .O(seg_15_18_sp4_r_v_b_17_62437)
  );
  Span4Mux_v4 t3473 (
    .I(seg_16_11_sp4_h_l_36_50315),
    .O(seg_16_15_sp4_v_b_1_61940)
  );
  Span4Mux_h4 t3474 (
    .I(seg_12_11_sp4_h_l_36_34991),
    .O(seg_16_11_sp4_h_l_36_50315)
  );
  LocalMux t3475 (
    .I(seg_20_6_sp4_v_b_12_76195),
    .O(seg_20_6_local_g1_4_79632)
  );
  Span4Mux_v1 t3476 (
    .I(seg_20_7_sp4_h_l_42_65153),
    .O(seg_20_6_sp4_v_b_12_76195)
  );
  Span4Mux_h4 t3477 (
    .I(seg_16_7_sp4_v_t_42_61454),
    .O(seg_20_7_sp4_h_l_42_65153)
  );
  Span4Mux_v4 t3478 (
    .I(seg_16_11_sp4_h_l_36_50315),
    .O(seg_16_7_sp4_v_t_42_61454)
  );
  LocalMux t3479 (
    .I(seg_20_7_sp4_h_r_7_79846),
    .O(seg_20_7_local_g0_7_79750)
  );
  CascadeMux t348 (
    .I(net_23706),
    .O(net_23706_cascademuxed)
  );
  Span4Mux_h0 t3480 (
    .I(seg_20_7_sp4_h_l_42_65153),
    .O(seg_20_7_sp4_h_r_7_79846)
  );
  LocalMux t3481 (
    .I(seg_8_14_sp4_v_b_16_31298),
    .O(seg_8_14_local_g1_0_35273)
  );
  Span4Mux_v3 t3482 (
    .I(seg_8_11_sp4_h_r_5_34997),
    .O(seg_8_14_sp4_v_b_16_31298)
  );
  LocalMux t3483 (
    .I(seg_2_7_sp4_r_v_b_10_11797),
    .O(seg_2_7_local_g2_2_12067)
  );
  Span4Mux_v1 t3484 (
    .I(seg_3_7_sp4_h_r_10_15976),
    .O(seg_2_7_sp4_r_v_b_10_11797)
  );
  Span4Mux_h4 t3485 (
    .I(seg_7_7_sp4_v_t_41_27438),
    .O(seg_3_7_sp4_h_r_10_15976)
  );
  Span4Mux_v4 t3486 (
    .I(seg_7_11_sp4_h_r_4_31165),
    .O(seg_7_7_sp4_v_t_41_27438)
  );
  LocalMux t3487 (
    .I(seg_3_6_sp4_v_b_23_11797),
    .O(seg_3_6_local_g1_7_15772)
  );
  Span4Mux_v1 t3488 (
    .I(seg_3_7_sp4_h_r_10_15976),
    .O(seg_3_6_sp4_v_b_23_11797)
  );
  LocalMux t3489 (
    .I(seg_3_18_sp4_v_b_17_13267),
    .O(seg_3_18_local_g0_1_17234)
  );
  CascadeMux t349 (
    .I(net_23736),
    .O(net_23736_cascademuxed)
  );
  Span4Mux_v3 t3490 (
    .I(seg_3_15_sp4_h_r_4_16964),
    .O(seg_3_18_sp4_v_b_17_13267)
  );
  Span4Mux_h4 t3491 (
    .I(seg_7_15_sp4_v_b_4_27846),
    .O(seg_3_15_sp4_h_r_4_16964)
  );
  Span4Mux_v4 t3492 (
    .I(seg_7_11_sp4_h_r_4_31165),
    .O(seg_7_15_sp4_v_b_4_27846)
  );
  LocalMux t3493 (
    .I(seg_4_7_sp4_h_r_23_15976),
    .O(seg_4_7_local_g1_7_19726)
  );
  Span4Mux_h3 t3494 (
    .I(seg_7_7_sp4_v_t_41_27438),
    .O(seg_4_7_sp4_h_r_23_15976)
  );
  LocalMux t3495 (
    .I(seg_7_5_sp4_v_b_24_27026),
    .O(seg_7_5_local_g2_0_30343)
  );
  Span4Mux_v2 t3496 (
    .I(seg_7_7_sp4_v_t_41_27438),
    .O(seg_7_5_sp4_v_b_24_27026)
  );
  LocalMux t3497 (
    .I(seg_7_15_sp4_v_b_4_27846),
    .O(seg_7_15_local_g0_4_31561)
  );
  LocalMux t3498 (
    .I(seg_7_15_sp4_v_b_4_27846),
    .O(seg_7_15_local_g1_4_31569)
  );
  LocalMux t3499 (
    .I(seg_15_6_sp4_v_b_14_57128),
    .O(seg_15_6_local_g0_6_61102)
  );
  CascadeMux t35 (
    .I(net_8155),
    .O(net_8155_cascademuxed)
  );
  CascadeMux t350 (
    .I(net_23964),
    .O(net_23964_cascademuxed)
  );
  Span4Mux_v1 t3500 (
    .I(seg_15_7_sp4_h_l_44_46002),
    .O(seg_15_6_sp4_v_b_14_57128)
  );
  Span4Mux_h4 t3501 (
    .I(seg_11_7_sp4_v_t_41_42300),
    .O(seg_15_7_sp4_h_l_44_46002)
  );
  Span4Mux_v4 t3502 (
    .I(seg_11_11_sp4_h_l_41_31165),
    .O(seg_11_7_sp4_v_t_41_42300)
  );
  LocalMux t3503 (
    .I(seg_3_6_sp4_v_b_12_11786),
    .O(seg_3_6_local_g0_4_15761)
  );
  Span4Mux_v1 t3504 (
    .I(seg_3_7_sp4_h_r_8_15984),
    .O(seg_3_6_sp4_v_b_12_11786)
  );
  Span4Mux_h4 t3505 (
    .I(seg_7_7_sp4_v_t_45_27442),
    .O(seg_3_7_sp4_h_r_8_15984)
  );
  Span4Mux_v4 t3506 (
    .I(seg_7_11_sp4_h_r_8_31169),
    .O(seg_7_7_sp4_v_t_45_27442)
  );
  LocalMux t3507 (
    .I(seg_7_5_sp4_v_b_28_27030),
    .O(seg_7_5_local_g3_4_30355)
  );
  Span4Mux_v2 t3508 (
    .I(seg_7_7_sp4_v_t_45_27442),
    .O(seg_7_5_sp4_v_b_28_27030)
  );
  LocalMux t3509 (
    .I(seg_5_14_sp4_r_v_b_20_24271),
    .O(seg_5_14_local_g3_4_24431)
  );
  CascadeMux t351 (
    .I(net_24081),
    .O(net_24081_cascademuxed)
  );
  Span4Mux_v3 t3510 (
    .I(seg_6_11_sp4_h_r_9_27738),
    .O(seg_5_14_sp4_r_v_b_20_24271)
  );
  LocalMux t3511 (
    .I(seg_10_4_sp4_v_b_36_37972),
    .O(seg_10_4_local_g3_4_41725)
  );
  Span4Mux_v3 t3512 (
    .I(seg_10_7_sp4_v_t_36_38464),
    .O(seg_10_4_sp4_v_b_36_37972)
  );
  LocalMux t3513 (
    .I(seg_12_7_sp4_h_r_25_42161),
    .O(seg_12_7_local_g2_1_49745)
  );
  Span4Mux_h2 t3514 (
    .I(seg_10_7_sp4_v_t_36_38464),
    .O(seg_12_7_sp4_h_r_25_42161)
  );
  LocalMux t3515 (
    .I(seg_13_6_sp4_r_v_b_18_53302),
    .O(seg_13_6_local_g3_2_53462)
  );
  Span4Mux_v1 t3516 (
    .I(seg_14_7_sp4_h_l_36_42161),
    .O(seg_13_6_sp4_r_v_b_18_53302)
  );
  Span4Mux_h4 t3517 (
    .I(seg_10_7_sp4_v_t_36_38464),
    .O(seg_14_7_sp4_h_l_36_42161)
  );
  LocalMux t3518 (
    .I(seg_13_7_sp4_h_r_36_42161),
    .O(seg_13_7_local_g2_4_53579)
  );
  Span4Mux_h3 t3519 (
    .I(seg_10_7_sp4_v_t_36_38464),
    .O(seg_13_7_sp4_h_r_36_42161)
  );
  CascadeMux t352 (
    .I(net_24087),
    .O(net_24087_cascademuxed)
  );
  LocalMux t3520 (
    .I(seg_13_7_sp4_h_r_36_42161),
    .O(seg_13_7_local_g3_4_53587)
  );
  LocalMux t3521 (
    .I(seg_14_5_sp4_v_b_30_53303),
    .O(seg_14_5_local_g2_6_57165)
  );
  Span4Mux_v2 t3522 (
    .I(seg_14_7_sp4_h_l_43_42168),
    .O(seg_14_5_sp4_v_b_30_53303)
  );
  Span4Mux_h4 t3523 (
    .I(seg_10_7_sp4_v_t_36_38464),
    .O(seg_14_7_sp4_h_l_43_42168)
  );
  LocalMux t3524 (
    .I(seg_14_5_sp4_v_b_31_53302),
    .O(seg_14_5_local_g2_7_57166)
  );
  Span4Mux_v2 t3525 (
    .I(seg_14_7_sp4_h_l_36_42161),
    .O(seg_14_5_sp4_v_b_31_53302)
  );
  LocalMux t3526 (
    .I(seg_14_5_sp4_v_b_31_53302),
    .O(seg_14_5_local_g3_7_57174)
  );
  LocalMux t3527 (
    .I(seg_14_6_sp4_v_b_18_53302),
    .O(seg_14_6_local_g1_2_57276)
  );
  Span4Mux_v1 t3528 (
    .I(seg_14_7_sp4_h_l_36_42161),
    .O(seg_14_6_sp4_v_b_18_53302)
  );
  LocalMux t3529 (
    .I(seg_14_6_sp4_v_b_19_53303),
    .O(seg_14_6_local_g1_3_57277)
  );
  CascadeMux t353 (
    .I(net_24216),
    .O(net_24216_cascademuxed)
  );
  Span4Mux_v1 t3530 (
    .I(seg_14_7_sp4_h_l_43_42168),
    .O(seg_14_6_sp4_v_b_19_53303)
  );
  LocalMux t3531 (
    .I(seg_2_8_sp4_h_r_0_12266),
    .O(seg_2_8_local_g0_0_12172)
  );
  Span4Mux_h4 t3532 (
    .I(seg_6_8_sp4_h_r_0_27421),
    .O(seg_2_8_sp4_h_r_0_12266)
  );
  Span4Mux_h4 t3533 (
    .I(seg_10_8_sp4_v_t_37_38588),
    .O(seg_6_8_sp4_h_r_0_27421)
  );
  LocalMux t3534 (
    .I(seg_2_8_sp4_h_r_0_12266),
    .O(seg_2_8_local_g1_0_12180)
  );
  LocalMux t3535 (
    .I(seg_2_8_sp4_h_r_3_12271),
    .O(seg_2_8_local_g1_3_12183)
  );
  Span4Mux_h4 t3536 (
    .I(seg_6_8_sp4_h_r_0_27421),
    .O(seg_2_8_sp4_h_r_3_12271)
  );
  LocalMux t3537 (
    .I(seg_10_4_sp4_h_r_5_41798),
    .O(seg_10_4_local_g1_5_41710)
  );
  Span4Mux_h0 t3538 (
    .I(seg_10_4_sp4_v_t_37_38096),
    .O(seg_10_4_sp4_h_r_5_41798)
  );
  Span4Mux_v4 t3539 (
    .I(seg_10_8_sp4_v_t_37_38588),
    .O(seg_10_4_sp4_v_t_37_38096)
  );
  CascadeMux t354 (
    .I(net_24333),
    .O(net_24333_cascademuxed)
  );
  LocalMux t3540 (
    .I(seg_10_19_sp4_v_b_17_39576),
    .O(seg_10_19_local_g1_1_43551)
  );
  Span4Mux_v3 t3541 (
    .I(seg_10_16_sp4_v_b_8_39088),
    .O(seg_10_19_sp4_v_b_17_39576)
  );
  Span4Mux_v4 t3542 (
    .I(seg_10_12_sp4_v_b_0_38588),
    .O(seg_10_16_sp4_v_b_8_39088)
  );
  LocalMux t3543 (
    .I(seg_12_4_sp4_h_r_29_41798),
    .O(seg_12_4_local_g2_5_49380)
  );
  Span4Mux_h2 t3544 (
    .I(seg_10_4_sp4_v_t_37_38096),
    .O(seg_12_4_sp4_h_r_29_41798)
  );
  LocalMux t3545 (
    .I(seg_12_4_sp4_h_r_29_41798),
    .O(seg_12_4_local_g3_5_49388)
  );
  LocalMux t3546 (
    .I(seg_13_7_sp4_r_v_b_13_53420),
    .O(seg_13_7_local_g2_5_53580)
  );
  Span4Mux_v1 t3547 (
    .I(seg_14_8_sp4_h_l_37_42283),
    .O(seg_13_7_sp4_r_v_b_13_53420)
  );
  Span4Mux_h4 t3548 (
    .I(seg_10_8_sp4_v_t_37_38588),
    .O(seg_14_8_sp4_h_l_37_42283)
  );
  LocalMux t3549 (
    .I(seg_13_7_sp4_r_v_b_19_53426),
    .O(seg_13_7_local_g3_3_53586)
  );
  CascadeMux t355 (
    .I(net_24438),
    .O(net_24438_cascademuxed)
  );
  Span4Mux_v1 t3550 (
    .I(seg_14_8_sp4_h_l_37_42283),
    .O(seg_13_7_sp4_r_v_b_19_53426)
  );
  LocalMux t3551 (
    .I(seg_14_5_sp4_v_b_43_53426),
    .O(seg_14_5_local_g2_3_57162)
  );
  Span4Mux_v3 t3552 (
    .I(seg_14_8_sp4_h_l_37_42283),
    .O(seg_14_5_sp4_v_b_43_53426)
  );
  LocalMux t3553 (
    .I(seg_14_5_sp4_v_b_37_53420),
    .O(seg_14_5_local_g3_5_57172)
  );
  Span4Mux_v3 t3554 (
    .I(seg_14_8_sp4_h_l_37_42283),
    .O(seg_14_5_sp4_v_b_37_53420)
  );
  LocalMux t3555 (
    .I(seg_14_6_sp4_v_b_30_53426),
    .O(seg_14_6_local_g2_6_57288)
  );
  Span4Mux_v2 t3556 (
    .I(seg_14_8_sp4_h_l_37_42283),
    .O(seg_14_6_sp4_v_b_30_53426)
  );
  LocalMux t3557 (
    .I(seg_14_6_sp4_v_b_30_53426),
    .O(seg_14_6_local_g3_6_57296)
  );
  LocalMux t3558 (
    .I(seg_2_8_sp4_h_r_1_12267),
    .O(seg_2_8_local_g1_1_12181)
  );
  Span4Mux_h4 t3559 (
    .I(seg_6_8_sp4_h_r_10_27423),
    .O(seg_2_8_sp4_h_r_1_12267)
  );
  CascadeMux t356 (
    .I(net_24462),
    .O(net_24462_cascademuxed)
  );
  Span4Mux_h4 t3560 (
    .I(seg_10_8_sp4_v_t_41_38592),
    .O(seg_6_8_sp4_h_r_10_27423)
  );
  LocalMux t3561 (
    .I(seg_12_4_sp4_h_r_33_41802),
    .O(seg_12_4_local_g3_1_49384)
  );
  Span4Mux_h2 t3562 (
    .I(seg_10_4_sp4_v_t_41_38100),
    .O(seg_12_4_sp4_h_r_33_41802)
  );
  Span4Mux_v4 t3563 (
    .I(seg_10_8_sp4_v_t_41_38592),
    .O(seg_10_4_sp4_v_t_41_38100)
  );
  LocalMux t3564 (
    .I(seg_2_7_sp4_h_r_20_7766),
    .O(seg_2_7_local_g0_4_12053)
  );
  Span4Mux_h3 t3565 (
    .I(seg_5_7_sp4_h_r_6_23644),
    .O(seg_2_7_sp4_h_r_20_7766)
  );
  Span4Mux_h4 t3566 (
    .I(seg_9_7_sp4_v_t_37_34634),
    .O(seg_5_7_sp4_h_r_6_23644)
  );
  LocalMux t3567 (
    .I(seg_4_6_sp4_r_v_b_19_19455),
    .O(seg_4_6_local_g3_3_19615)
  );
  Span4Mux_v1 t3568 (
    .I(seg_5_7_sp4_h_r_6_23644),
    .O(seg_4_6_sp4_r_v_b_19_19455)
  );
  LocalMux t3569 (
    .I(seg_5_3_sp4_h_r_11_23147),
    .O(seg_5_3_local_g1_3_23061)
  );
  CascadeMux t357 (
    .I(net_24696),
    .O(net_24696_cascademuxed)
  );
  Span4Mux_h0 t3570 (
    .I(seg_5_3_sp4_v_t_43_19455),
    .O(seg_5_3_sp4_h_r_11_23147)
  );
  Span4Mux_v4 t3571 (
    .I(seg_5_7_sp4_h_r_6_23644),
    .O(seg_5_3_sp4_v_t_43_19455)
  );
  LocalMux t3572 (
    .I(seg_5_7_sp4_h_r_6_23644),
    .O(seg_5_7_local_g0_6_23548)
  );
  LocalMux t3573 (
    .I(seg_5_7_sp4_h_r_6_23644),
    .O(seg_5_7_local_g1_6_23556)
  );
  LocalMux t3574 (
    .I(seg_5_14_sp4_v_b_13_20433),
    .O(seg_5_14_local_g1_5_24416)
  );
  Span4Mux_v3 t3575 (
    .I(seg_5_11_sp4_h_r_0_24128),
    .O(seg_5_14_sp4_v_b_13_20433)
  );
  Span4Mux_h4 t3576 (
    .I(seg_9_11_sp4_v_b_0_34634),
    .O(seg_5_11_sp4_h_r_0_24128)
  );
  LocalMux t3577 (
    .I(seg_8_3_sp4_r_v_b_11_33765),
    .O(seg_8_3_local_g2_3_33931)
  );
  Span4Mux_v1 t3578 (
    .I(seg_9_3_sp4_v_t_45_34150),
    .O(seg_8_3_sp4_r_v_b_11_33765)
  );
  Span4Mux_v4 t3579 (
    .I(seg_9_7_sp4_v_t_37_34634),
    .O(seg_9_3_sp4_v_t_45_34150)
  );
  CascadeMux t358 (
    .I(net_24714),
    .O(net_24714_cascademuxed)
  );
  LocalMux t3580 (
    .I(seg_9_3_sp4_h_r_8_37847),
    .O(seg_9_3_local_g0_0_37743)
  );
  Span4Mux_h0 t3581 (
    .I(seg_9_3_sp4_v_t_45_34150),
    .O(seg_9_3_sp4_h_r_8_37847)
  );
  LocalMux t3582 (
    .I(seg_9_4_sp4_v_b_45_34150),
    .O(seg_9_4_local_g3_5_37895)
  );
  Span4Mux_v3 t3583 (
    .I(seg_9_7_sp4_v_t_37_34634),
    .O(seg_9_4_sp4_v_b_45_34150)
  );
  LocalMux t3584 (
    .I(seg_4_5_sp4_r_v_b_36_19571),
    .O(seg_4_5_local_g2_4_19485)
  );
  Span4Mux_v3 t3585 (
    .I(seg_5_8_sp4_h_r_1_23760),
    .O(seg_4_5_sp4_r_v_b_36_19571)
  );
  Span4Mux_h4 t3586 (
    .I(seg_9_8_sp4_v_t_36_34756),
    .O(seg_5_8_sp4_h_r_1_23760)
  );
  LocalMux t3587 (
    .I(seg_4_6_sp4_r_v_b_24_19572),
    .O(seg_4_6_local_g0_0_19588)
  );
  Span4Mux_v2 t3588 (
    .I(seg_5_8_sp4_h_r_7_23768),
    .O(seg_4_6_sp4_r_v_b_24_19572)
  );
  Span4Mux_h4 t3589 (
    .I(seg_9_8_sp4_v_t_36_34756),
    .O(seg_5_8_sp4_h_r_7_23768)
  );
  CascadeMux t359 (
    .I(net_24720),
    .O(net_24720_cascademuxed)
  );
  LocalMux t3590 (
    .I(seg_4_7_sp4_r_v_b_18_19577),
    .O(seg_4_7_local_g3_2_19737)
  );
  Span4Mux_v1 t3591 (
    .I(seg_5_8_sp4_h_r_7_23768),
    .O(seg_4_7_sp4_r_v_b_18_19577)
  );
  LocalMux t3592 (
    .I(seg_5_3_sp4_v_b_21_19083),
    .O(seg_5_3_local_g1_5_23063)
  );
  Span4Mux_v1 t3593 (
    .I(seg_5_4_sp4_v_t_37_19572),
    .O(seg_5_3_sp4_v_b_21_19083)
  );
  Span4Mux_v4 t3594 (
    .I(seg_5_8_sp4_h_r_7_23768),
    .O(seg_5_4_sp4_v_t_37_19572)
  );
  LocalMux t3595 (
    .I(seg_5_7_sp4_v_b_13_19572),
    .O(seg_5_7_local_g0_5_23547)
  );
  Span4Mux_v1 t3596 (
    .I(seg_5_8_sp4_h_r_7_23768),
    .O(seg_5_7_sp4_v_b_13_19572)
  );
  LocalMux t3597 (
    .I(seg_5_16_sp4_v_b_0_20556),
    .O(seg_5_16_local_g1_0_24657)
  );
  Span4Mux_v4 t3598 (
    .I(seg_5_12_sp4_h_r_6_24259),
    .O(seg_5_16_sp4_v_b_0_20556)
  );
  Span4Mux_h4 t3599 (
    .I(seg_9_12_sp4_v_b_1_34756),
    .O(seg_5_12_sp4_h_r_6_24259)
  );
  CascadeMux t360 (
    .I(net_24726),
    .O(net_24726_cascademuxed)
  );
  LocalMux t3600 (
    .I(seg_5_16_sp4_v_b_1_20555),
    .O(seg_5_16_local_g1_1_24658)
  );
  Span4Mux_v4 t3601 (
    .I(seg_5_12_sp4_h_r_1_24252),
    .O(seg_5_16_sp4_v_b_1_20555)
  );
  Span4Mux_h4 t3602 (
    .I(seg_9_12_sp4_v_b_1_34756),
    .O(seg_5_12_sp4_h_r_1_24252)
  );
  LocalMux t3603 (
    .I(seg_8_3_sp4_r_v_b_17_33772),
    .O(seg_8_3_local_g3_1_33937)
  );
  Span4Mux_v1 t3604 (
    .I(seg_9_4_sp4_v_t_36_34264),
    .O(seg_8_3_sp4_r_v_b_17_33772)
  );
  Span4Mux_v4 t3605 (
    .I(seg_9_8_sp4_v_t_36_34756),
    .O(seg_9_4_sp4_v_t_36_34264)
  );
  LocalMux t3606 (
    .I(seg_8_16_sp4_r_v_b_9_35256),
    .O(seg_8_16_local_g2_1_35528)
  );
  Span4Mux_v4 t3607 (
    .I(seg_9_12_sp4_v_b_1_34756),
    .O(seg_8_16_sp4_r_v_b_9_35256)
  );
  LocalMux t3608 (
    .I(seg_9_3_sp4_v_b_17_33772),
    .O(seg_9_3_local_g1_1_37752)
  );
  Span4Mux_v1 t3609 (
    .I(seg_9_4_sp4_v_t_36_34264),
    .O(seg_9_3_sp4_v_b_17_33772)
  );
  CascadeMux t361 (
    .I(net_24813),
    .O(net_24813_cascademuxed)
  );
  LocalMux t3610 (
    .I(seg_9_4_sp4_h_r_6_37968),
    .O(seg_9_4_local_g1_6_37880)
  );
  Span4Mux_h0 t3611 (
    .I(seg_9_4_sp4_v_t_36_34264),
    .O(seg_9_4_sp4_h_r_6_37968)
  );
  LocalMux t3612 (
    .I(seg_10_4_sp4_h_r_19_37968),
    .O(seg_10_4_local_g1_3_41708)
  );
  Span4Mux_h1 t3613 (
    .I(seg_9_4_sp4_v_t_36_34264),
    .O(seg_10_4_sp4_h_r_19_37968)
  );
  LocalMux t3614 (
    .I(seg_12_7_sp4_r_v_b_19_49595),
    .O(seg_12_7_local_g3_3_49755)
  );
  Span4Mux_v1 t3615 (
    .I(seg_13_8_sp4_h_l_43_38460),
    .O(seg_12_7_sp4_r_v_b_19_49595)
  );
  Span4Mux_h4 t3616 (
    .I(seg_9_8_sp4_v_t_36_34756),
    .O(seg_13_8_sp4_h_l_43_38460)
  );
  LocalMux t3617 (
    .I(seg_13_6_sp4_v_b_30_49595),
    .O(seg_13_6_local_g2_6_53458)
  );
  Span4Mux_v2 t3618 (
    .I(seg_13_8_sp4_h_l_43_38460),
    .O(seg_13_6_sp4_v_b_30_49595)
  );
  LocalMux t3619 (
    .I(seg_2_8_sp4_h_r_18_7911),
    .O(seg_2_8_local_g1_2_12182)
  );
  CascadeMux t362 (
    .I(net_24948),
    .O(net_24948_cascademuxed)
  );
  Span4Mux_h3 t3620 (
    .I(seg_5_8_sp4_h_r_11_23762),
    .O(seg_2_8_sp4_h_r_18_7911)
  );
  Span4Mux_h4 t3621 (
    .I(seg_9_8_sp4_v_t_40_34760),
    .O(seg_5_8_sp4_h_r_11_23762)
  );
  LocalMux t3622 (
    .I(seg_4_5_sp4_r_v_b_46_19581),
    .O(seg_4_5_local_g3_6_19495)
  );
  Span4Mux_v3 t3623 (
    .I(seg_5_8_sp4_h_r_11_23762),
    .O(seg_4_5_sp4_r_v_b_46_19581)
  );
  LocalMux t3624 (
    .I(seg_4_7_sp4_r_v_b_17_19576),
    .O(seg_4_7_local_g3_1_19736)
  );
  Span4Mux_v1 t3625 (
    .I(seg_5_8_sp4_h_r_11_23762),
    .O(seg_4_7_sp4_r_v_b_17_19576)
  );
  LocalMux t3626 (
    .I(seg_8_16_sp4_r_v_b_17_35376),
    .O(seg_8_16_local_g3_1_35536)
  );
  Span4Mux_v3 t3627 (
    .I(seg_9_13_sp4_v_b_4_34884),
    .O(seg_8_16_sp4_r_v_b_17_35376)
  );
  LocalMux t3628 (
    .I(seg_4_18_sp4_r_v_b_3_20803),
    .O(seg_4_18_local_g1_3_21075)
  );
  Span4Mux_v4 t3629 (
    .I(seg_5_14_sp4_h_r_9_24508),
    .O(seg_4_18_sp4_r_v_b_3_20803)
  );
  CascadeMux t363 (
    .I(net_25053),
    .O(net_25053_cascademuxed)
  );
  Span4Mux_h4 t3630 (
    .I(seg_9_14_sp4_v_b_9_35010),
    .O(seg_5_14_sp4_h_r_9_24508)
  );
  LocalMux t3631 (
    .I(seg_8_14_sp4_r_v_b_9_35010),
    .O(seg_8_14_local_g2_1_35282)
  );
  LocalMux t3632 (
    .I(seg_8_12_neigh_op_rgt_5_34983),
    .O(seg_8_12_local_g2_5_35040)
  );
  LocalMux t3633 (
    .I(seg_8_15_sp4_v_b_22_31427),
    .O(seg_8_15_local_g0_6_35394)
  );
  Span4Mux_v3 t3634 (
    .I(seg_8_12_sp4_h_r_5_35120),
    .O(seg_8_15_sp4_v_b_22_31427)
  );
  LocalMux t3635 (
    .I(seg_8_15_sp4_v_b_18_31423),
    .O(seg_8_15_local_g0_2_35390)
  );
  Span4Mux_v3 t3636 (
    .I(seg_8_12_sp4_h_r_7_35122),
    .O(seg_8_15_sp4_v_b_18_31423)
  );
  LocalMux t3637 (
    .I(seg_8_15_sp4_r_v_b_5_35129),
    .O(seg_8_15_local_g1_5_35401)
  );
  LocalMux t3638 (
    .I(seg_9_13_lutff_3_out_35104),
    .O(seg_9_13_local_g3_3_39000)
  );
  LocalMux t3639 (
    .I(seg_11_13_sp4_h_r_34_39069),
    .O(seg_11_13_local_g3_2_46661)
  );
  CascadeMux t364 (
    .I(net_25077),
    .O(net_25077_cascademuxed)
  );
  LocalMux t3640 (
    .I(seg_8_15_sp4_r_v_b_4_35130),
    .O(seg_8_15_local_g1_4_35400)
  );
  LocalMux t3641 (
    .I(seg_8_15_neigh_op_bnr_0_35224),
    .O(seg_8_15_local_g1_0_35396)
  );
  LocalMux t3642 (
    .I(seg_10_15_neigh_op_bnl_2_35226),
    .O(seg_10_15_local_g3_2_43076)
  );
  LocalMux t3643 (
    .I(seg_9_14_lutff_3_out_35227),
    .O(seg_9_14_local_g2_3_39115)
  );
  LocalMux t3644 (
    .I(seg_9_15_neigh_op_bot_4_35228),
    .O(seg_9_15_local_g1_4_39231)
  );
  LocalMux t3645 (
    .I(seg_9_15_neigh_op_bot_7_35231),
    .O(seg_9_15_local_g1_7_39234)
  );
  LocalMux t3646 (
    .I(seg_11_15_sp4_v_b_39_43159),
    .O(seg_11_15_local_g2_7_46904)
  );
  Span4Mux_v1 t3647 (
    .I(seg_11_14_sp4_h_l_39_31532),
    .O(seg_11_15_sp4_v_b_39_43159)
  );
  LocalMux t3648 (
    .I(seg_8_15_neigh_op_rgt_0_35347),
    .O(seg_8_15_local_g2_0_35404)
  );
  LocalMux t3649 (
    .I(seg_8_15_neigh_op_rgt_1_35348),
    .O(seg_8_15_local_g2_1_35405)
  );
  CascadeMux t365 (
    .I(net_26885),
    .O(net_26885_cascademuxed)
  );
  LocalMux t3650 (
    .I(seg_8_15_neigh_op_rgt_3_35350),
    .O(seg_8_15_local_g3_3_35415)
  );
  LocalMux t3651 (
    .I(seg_8_15_neigh_op_rgt_4_35351),
    .O(seg_8_15_local_g3_4_35416)
  );
  LocalMux t3652 (
    .I(seg_8_15_neigh_op_rgt_5_35352),
    .O(seg_8_15_local_g3_5_35417)
  );
  LocalMux t3653 (
    .I(seg_8_15_neigh_op_rgt_6_35353),
    .O(seg_8_15_local_g2_6_35410)
  );
  LocalMux t3654 (
    .I(seg_8_15_neigh_op_rgt_7_35354),
    .O(seg_8_15_local_g3_7_35419)
  );
  LocalMux t3655 (
    .I(seg_9_18_sp4_r_v_b_12_39448),
    .O(seg_9_18_local_g2_4_39608)
  );
  Span4Mux_v3 t3656 (
    .I(seg_10_15_sp4_h_l_36_28136),
    .O(seg_9_18_sp4_r_v_b_12_39448)
  );
  LocalMux t3657 (
    .I(seg_9_18_sp4_v_b_24_35741),
    .O(seg_9_18_local_g2_0_39604)
  );
  Span4Mux_v2 t3658 (
    .I(seg_9_16_sp4_h_r_0_39436),
    .O(seg_9_18_sp4_v_b_24_35741)
  );
  LocalMux t3659 (
    .I(seg_9_18_sp4_r_v_b_7_39331),
    .O(seg_9_18_local_g1_7_39603)
  );
  CascadeMux t366 (
    .I(net_26886),
    .O(net_26886_cascademuxed)
  );
  LocalMux t3660 (
    .I(seg_9_18_sp4_r_v_b_17_39453),
    .O(seg_9_18_local_g3_1_39613)
  );
  LocalMux t3661 (
    .I(seg_9_18_sp4_r_v_b_19_39455),
    .O(seg_9_18_local_g3_3_39615)
  );
  LocalMux t3662 (
    .I(seg_9_18_sp4_v_b_14_35619),
    .O(seg_9_18_local_g0_6_39594)
  );
  LocalMux t3663 (
    .I(seg_9_17_lutff_0_out_35593),
    .O(seg_9_17_local_g2_0_39481)
  );
  LocalMux t3664 (
    .I(seg_9_18_neigh_op_bot_2_35595),
    .O(seg_9_18_local_g1_2_39598)
  );
  LocalMux t3665 (
    .I(seg_9_17_lutff_3_out_35596),
    .O(seg_9_17_local_g3_3_39492)
  );
  LocalMux t3666 (
    .I(seg_9_18_sp4_r_v_b_22_39458),
    .O(seg_9_18_local_g3_6_39618)
  );
  LocalMux t3667 (
    .I(seg_10_18_neigh_op_lft_0_35716),
    .O(seg_10_18_local_g0_0_43419)
  );
  LocalMux t3668 (
    .I(seg_10_18_neigh_op_lft_2_35718),
    .O(seg_10_18_local_g0_2_43421)
  );
  LocalMux t3669 (
    .I(seg_10_18_neigh_op_lft_5_35721),
    .O(seg_10_18_local_g1_5_43432)
  );
  CascadeMux t367 (
    .I(net_26888),
    .O(net_26888_cascademuxed)
  );
  LocalMux t3670 (
    .I(seg_10_18_neigh_op_lft_6_35722),
    .O(seg_10_18_local_g0_6_43425)
  );
  LocalMux t3671 (
    .I(seg_10_18_neigh_op_lft_7_35723),
    .O(seg_10_18_local_g1_7_43434)
  );
  LocalMux t3672 (
    .I(seg_11_16_sp4_h_r_17_43273),
    .O(seg_11_16_local_g1_1_47013)
  );
  Span4Mux_h1 t3673 (
    .I(seg_10_16_sp4_v_t_46_39581),
    .O(seg_11_16_sp4_h_r_17_43273)
  );
  LocalMux t3674 (
    .I(seg_11_2_neigh_op_bnl_1_37416),
    .O(seg_11_2_local_g2_1_45299)
  );
  LocalMux t3675 (
    .I(seg_11_2_neigh_op_bnl_2_37417),
    .O(seg_11_2_local_g3_2_45308)
  );
  LocalMux t3676 (
    .I(seg_10_1_lutff_5_out_37420),
    .O(seg_10_1_local_g2_5_41309)
  );
  LocalMux t3677 (
    .I(seg_10_1_lutff_6_out_37421),
    .O(seg_10_1_local_g0_6_41294)
  );
  LocalMux t3678 (
    .I(seg_11_2_neigh_op_bnl_7_37422),
    .O(seg_11_2_local_g2_7_45305)
  );
  LocalMux t3679 (
    .I(seg_13_4_sp4_h_r_28_45628),
    .O(seg_13_4_local_g2_4_53210)
  );
  CascadeMux t368 (
    .I(net_26889),
    .O(net_26889_cascademuxed)
  );
  Span4Mux_h2 t3680 (
    .I(seg_11_4_sp4_v_b_10_41440),
    .O(seg_13_4_sp4_h_r_28_45628)
  );
  LocalMux t3681 (
    .I(seg_10_2_lutff_0_out_37543),
    .O(seg_10_2_local_g3_0_41475)
  );
  LocalMux t3682 (
    .I(seg_11_3_neigh_op_bnl_1_37544),
    .O(seg_11_3_local_g3_1_45430)
  );
  LocalMux t3683 (
    .I(seg_10_2_lutff_2_out_37545),
    .O(seg_10_2_local_g3_2_41477)
  );
  LocalMux t3684 (
    .I(seg_10_2_lutff_3_out_37546),
    .O(seg_10_2_local_g2_3_41470)
  );
  LocalMux t3685 (
    .I(seg_11_3_neigh_op_bnl_4_37547),
    .O(seg_11_3_local_g2_4_45425)
  );
  LocalMux t3686 (
    .I(seg_10_1_neigh_op_top_5_37548),
    .O(seg_10_1_local_g0_5_41293)
  );
  LocalMux t3687 (
    .I(seg_10_2_lutff_6_out_37549),
    .O(seg_10_2_local_g0_6_41457)
  );
  LocalMux t3688 (
    .I(seg_10_1_neigh_op_top_7_37550),
    .O(seg_10_1_local_g1_7_41303)
  );
  LocalMux t3689 (
    .I(seg_11_3_neigh_op_lft_0_37702),
    .O(seg_11_3_local_g1_0_45413)
  );
  CascadeMux t369 (
    .I(net_26890),
    .O(net_26890_cascademuxed)
  );
  LocalMux t3690 (
    .I(seg_11_3_neigh_op_lft_1_37703),
    .O(seg_11_3_local_g1_1_45414)
  );
  LocalMux t3691 (
    .I(seg_11_3_neigh_op_lft_2_37704),
    .O(seg_11_3_local_g1_2_45415)
  );
  LocalMux t3692 (
    .I(seg_11_3_neigh_op_lft_3_37705),
    .O(seg_11_3_local_g0_3_45408)
  );
  LocalMux t3693 (
    .I(seg_11_3_neigh_op_lft_4_37706),
    .O(seg_11_3_local_g1_4_45417)
  );
  LocalMux t3694 (
    .I(seg_11_3_neigh_op_lft_5_37707),
    .O(seg_11_3_local_g1_5_45418)
  );
  LocalMux t3695 (
    .I(seg_11_3_neigh_op_lft_6_37708),
    .O(seg_11_3_local_g0_6_45411)
  );
  LocalMux t3696 (
    .I(seg_11_3_neigh_op_lft_7_37709),
    .O(seg_11_3_local_g1_7_45420)
  );
  LocalMux t3697 (
    .I(seg_12_4_sp4_h_r_31_41800),
    .O(seg_12_4_local_g3_7_49390)
  );
  Span4Mux_h2 t3698 (
    .I(seg_10_4_sp4_v_b_1_37597),
    .O(seg_12_4_sp4_h_r_31_41800)
  );
  LocalMux t3699 (
    .I(seg_10_4_lutff_1_out_37826),
    .O(seg_10_4_local_g2_1_41714)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t37 (
    .carryinitin(),
    .carryinitout(t36)
  );
  CascadeMux t370 (
    .I(net_26891),
    .O(net_26891_cascademuxed)
  );
  LocalMux t3700 (
    .I(seg_9_4_neigh_op_rgt_3_37828),
    .O(seg_9_4_local_g2_3_37885)
  );
  LocalMux t3701 (
    .I(seg_10_4_lutff_6_out_37831),
    .O(seg_10_4_local_g3_6_41727)
  );
  LocalMux t3702 (
    .I(seg_10_19_sp12_v_b_11_42774),
    .O(seg_10_19_local_g3_3_43569)
  );
  Span12Mux_v7 t3703 (
    .I(seg_10_12_sp12_v_b_0_41270),
    .O(seg_10_19_sp12_v_b_11_42774)
  );
  LocalMux t3704 (
    .I(seg_12_4_sp4_h_r_34_41793),
    .O(seg_12_4_local_g3_2_49385)
  );
  LocalMux t3705 (
    .I(seg_15_6_sp4_h_r_10_61192),
    .O(seg_15_6_local_g1_2_61106)
  );
  Span4Mux_h0 t3706 (
    .I(seg_15_6_sp4_h_l_42_45877),
    .O(seg_15_6_sp4_h_r_10_61192)
  );
  Span4Mux_h4 t3707 (
    .I(seg_11_6_sp4_v_b_7_41686),
    .O(seg_15_6_sp4_h_l_42_45877)
  );
  LocalMux t3708 (
    .I(seg_10_5_lutff_4_out_37952),
    .O(seg_10_5_local_g1_4_41832)
  );
  LocalMux t3709 (
    .I(seg_10_5_lutff_5_out_37953),
    .O(seg_10_5_local_g3_5_41849)
  );
  LocalMux t3710 (
    .I(seg_11_5_neigh_op_lft_7_37955),
    .O(seg_11_5_local_g0_7_45658)
  );
  LocalMux t3711 (
    .I(seg_10_3_sp4_v_b_36_37849),
    .O(seg_10_3_local_g2_4_41594)
  );
  LocalMux t3712 (
    .I(seg_10_2_sp4_v_b_39_37729),
    .O(seg_10_2_local_g2_7_41474)
  );
  LocalMux t3713 (
    .I(seg_15_6_sp4_h_r_16_57367),
    .O(seg_15_6_local_g0_0_61096)
  );
  Span4Mux_h1 t3714 (
    .I(seg_14_6_sp4_h_l_39_42041),
    .O(seg_15_6_sp4_h_r_16_57367)
  );
  LocalMux t3715 (
    .I(seg_15_6_sp4_h_r_45_49709),
    .O(seg_15_6_local_g2_5_61117)
  );
  Span4Mux_h3 t3716 (
    .I(seg_12_6_sp4_h_l_37_34375),
    .O(seg_15_6_sp4_h_r_45_49709)
  );
  LocalMux t3717 (
    .I(seg_10_19_sp4_v_b_15_39574),
    .O(seg_10_19_local_g0_7_43549)
  );
  Span4Mux_v3 t3718 (
    .I(seg_10_16_sp4_v_b_2_39082),
    .O(seg_10_19_sp4_v_b_15_39574)
  );
  Span4Mux_v4 t3719 (
    .I(seg_10_12_sp4_v_b_6_38594),
    .O(seg_10_16_sp4_v_b_2_39082)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t372 (
    .carryinitin(),
    .carryinitout(t371)
  );
  Span4Mux_v4 t3720 (
    .I(seg_10_8_sp4_v_b_6_38102),
    .O(seg_10_12_sp4_v_b_6_38594)
  );
  LocalMux t3721 (
    .I(seg_11_7_neigh_op_lft_0_38194),
    .O(seg_11_7_local_g1_0_45905)
  );
  LocalMux t3722 (
    .I(seg_11_6_neigh_op_tnl_1_38195),
    .O(seg_11_6_local_g2_1_45791)
  );
  LocalMux t3723 (
    .I(seg_11_6_neigh_op_tnl_3_38197),
    .O(seg_11_6_local_g2_3_45793)
  );
  LocalMux t3724 (
    .I(seg_10_7_lutff_7_out_38201),
    .O(seg_10_7_local_g0_7_42073)
  );
  LocalMux t3725 (
    .I(seg_12_7_sp4_h_r_40_38336),
    .O(seg_12_7_local_g3_0_49752)
  );
  LocalMux t3726 (
    .I(seg_13_5_sp4_v_b_35_49475),
    .O(seg_13_5_local_g2_3_53332)
  );
  Span4Mux_v2 t3727 (
    .I(seg_13_7_sp4_h_l_40_38336),
    .O(seg_13_5_sp4_v_b_35_49475)
  );
  LocalMux t3728 (
    .I(seg_13_6_sp4_v_b_22_49475),
    .O(seg_13_6_local_g1_6_53450)
  );
  Span4Mux_v1 t3729 (
    .I(seg_13_7_sp4_h_l_40_38336),
    .O(seg_13_6_sp4_v_b_22_49475)
  );
  CascadeMux t373 (
    .I(net_26987),
    .O(net_26987_cascademuxed)
  );
  LocalMux t3730 (
    .I(seg_0_12_sp4_v_b_42_2510),
    .O(seg_0_12_local_g3_2_2546)
  );
  Span4Mux_v1 t3731 (
    .I(seg_0_11_sp4_v_b_4_1657),
    .O(seg_0_12_sp4_v_b_42_2510)
  );
  Span4Mux_v4 t3732 (
    .I(seg_0_7_sp4_h_r_4_1626),
    .O(seg_0_11_sp4_v_b_4_1657)
  );
  Span4Mux_h4 t3733 (
    .I(seg_4_7_sp4_h_r_8_19815),
    .O(seg_0_7_sp4_h_r_4_1626)
  );
  Span4Mux_h4 t3734 (
    .I(seg_8_7_sp4_h_r_0_34498),
    .O(seg_4_7_sp4_h_r_8_19815)
  );
  LocalMux t3735 (
    .I(seg_15_5_sp4_h_r_2_61071),
    .O(seg_15_5_local_g1_2_60983)
  );
  Span4Mux_h0 t3736 (
    .I(seg_15_5_sp4_h_l_39_45749),
    .O(seg_15_5_sp4_h_r_2_61071)
  );
  Span4Mux_h4 t3737 (
    .I(seg_11_5_sp4_v_t_44_42057),
    .O(seg_15_5_sp4_h_l_39_45749)
  );
  LocalMux t3738 (
    .I(seg_10_2_sp4_v_b_23_37595),
    .O(seg_10_2_local_g0_7_41458)
  );
  Span4Mux_v1 t3739 (
    .I(seg_10_3_sp4_v_t_47_37983),
    .O(seg_10_2_sp4_v_b_23_37595)
  );
  CascadeMux t374 (
    .I(net_26988),
    .O(net_26988_cascademuxed)
  );
  LocalMux t3740 (
    .I(seg_0_25_sp4_h_r_24_5470),
    .O(seg_0_25_local_g3_0_5345)
  );
  Span4Mux_h2 t3741 (
    .I(seg_2_25_sp4_h_r_9_14368),
    .O(seg_0_25_sp4_h_r_24_5470)
  );
  Span4Mux_h4 t3742 (
    .I(seg_6_25_sp4_h_r_1_29156),
    .O(seg_2_25_sp4_h_r_9_14368)
  );
  Span4Mux_h4 t3743 (
    .I(seg_10_25_sp4_v_b_8_40195),
    .O(seg_6_25_sp4_h_r_1_29156)
  );
  Span4Mux_v4 t3744 (
    .I(seg_10_21_sp4_v_b_0_39695),
    .O(seg_10_25_sp4_v_b_8_40195)
  );
  Span4Mux_v4 t3745 (
    .I(seg_10_17_sp4_v_b_0_39203),
    .O(seg_10_21_sp4_v_b_0_39695)
  );
  Span4Mux_v4 t3746 (
    .I(seg_10_13_sp4_v_b_0_38711),
    .O(seg_10_17_sp4_v_b_0_39203)
  );
  Span4Mux_v4 t3747 (
    .I(seg_10_9_sp4_v_b_0_38219),
    .O(seg_10_13_sp4_v_b_0_38711)
  );
  LocalMux t3748 (
    .I(seg_10_8_lutff_1_out_38318),
    .O(seg_10_8_local_g1_1_42198)
  );
  LocalMux t3749 (
    .I(seg_11_8_neigh_op_lft_3_38320),
    .O(seg_11_8_local_g1_3_46031)
  );
  CascadeMux t375 (
    .I(net_26990),
    .O(net_26990_cascademuxed)
  );
  LocalMux t3750 (
    .I(seg_10_7_neigh_op_top_4_38321),
    .O(seg_10_7_local_g0_4_42070)
  );
  LocalMux t3751 (
    .I(seg_10_8_lutff_5_out_38322),
    .O(seg_10_8_local_g3_5_42218)
  );
  LocalMux t3752 (
    .I(seg_11_8_neigh_op_lft_6_38323),
    .O(seg_11_8_local_g1_6_46034)
  );
  LocalMux t3753 (
    .I(seg_10_9_neigh_op_bot_7_38324),
    .O(seg_10_9_local_g0_7_42319)
  );
  LocalMux t3754 (
    .I(seg_12_7_sp4_r_v_b_14_49590),
    .O(seg_12_7_local_g2_6_49750)
  );
  Span4Mux_v1 t3755 (
    .I(seg_13_8_sp4_h_l_38_38457),
    .O(seg_12_7_sp4_r_v_b_14_49590)
  );
  LocalMux t3756 (
    .I(seg_13_3_sp4_v_b_22_49101),
    .O(seg_13_3_local_g0_6_53073)
  );
  Span4Mux_v1 t3757 (
    .I(seg_13_4_sp4_v_t_38_49590),
    .O(seg_13_3_sp4_v_b_22_49101)
  );
  Span4Mux_v4 t3758 (
    .I(seg_13_8_sp4_h_l_38_38457),
    .O(seg_13_4_sp4_v_t_38_49590)
  );
  LocalMux t3759 (
    .I(seg_12_4_sp4_h_r_23_45624),
    .O(seg_12_4_local_g0_7_49366)
  );
  CascadeMux t376 (
    .I(net_26991),
    .O(net_26991_cascademuxed)
  );
  Span4Mux_h1 t3760 (
    .I(seg_11_4_sp4_v_t_40_41930),
    .O(seg_12_4_sp4_h_r_23_45624)
  );
  Span4Mux_v4 t3761 (
    .I(seg_11_8_sp4_h_l_46_30793),
    .O(seg_11_4_sp4_v_t_40_41930)
  );
  LocalMux t3762 (
    .I(seg_11_4_sp4_h_r_6_45630),
    .O(seg_11_4_local_g0_6_45534)
  );
  Span4Mux_h0 t3763 (
    .I(seg_11_4_sp4_v_t_36_41926),
    .O(seg_11_4_sp4_h_r_6_45630)
  );
  LocalMux t3764 (
    .I(seg_11_19_sp4_v_b_9_43287),
    .O(seg_11_19_local_g1_1_47382)
  );
  Span4Mux_v4 t3765 (
    .I(seg_11_15_sp4_v_b_1_42787),
    .O(seg_11_19_sp4_v_b_9_43287)
  );
  Span4Mux_v4 t3766 (
    .I(seg_11_11_sp4_v_b_10_42306),
    .O(seg_11_15_sp4_v_b_1_42787)
  );
  LocalMux t3767 (
    .I(seg_10_19_sp12_v_b_2_42281),
    .O(seg_10_19_local_g3_2_43568)
  );
  LocalMux t3768 (
    .I(seg_10_10_lutff_1_out_38564),
    .O(seg_10_10_local_g0_1_42436)
  );
  LocalMux t3769 (
    .I(seg_10_10_lutff_3_out_38566),
    .O(seg_10_10_local_g2_3_42454)
  );
  CascadeMux t377 (
    .I(net_26992),
    .O(net_26992_cascademuxed)
  );
  LocalMux t3770 (
    .I(seg_10_10_lutff_5_out_38568),
    .O(seg_10_10_local_g2_5_42456)
  );
  LocalMux t3771 (
    .I(seg_0_25_sp12_v_b_19_4816),
    .O(seg_0_25_local_g2_3_5340)
  );
  Span12Mux_v3 t3772 (
    .I(seg_0_22_sp12_v_b_0_2225),
    .O(seg_0_25_sp12_v_b_19_4816)
  );
  Span12Mux_v12 t3773 (
    .I(seg_0_10_sp12_h_r_0_2200),
    .O(seg_0_22_sp12_v_b_0_2225)
  );
  LocalMux t3774 (
    .I(seg_9_14_sp4_r_v_b_6_38840),
    .O(seg_9_14_local_g1_6_39110)
  );
  Span4Mux_v4 t3775 (
    .I(seg_10_10_sp4_h_r_0_42529),
    .O(seg_9_14_sp4_r_v_b_6_38840)
  );
  LocalMux t3776 (
    .I(seg_9_14_sp4_v_b_3_35004),
    .O(seg_9_14_local_g0_3_39099)
  );
  Span4Mux_v4 t3777 (
    .I(seg_9_10_sp4_h_r_3_38703),
    .O(seg_9_14_sp4_v_b_3_35004)
  );
  LocalMux t3778 (
    .I(seg_0_12_sp4_v_b_24_2299),
    .O(seg_0_12_local_g3_0_2544)
  );
  Span4Mux_v2 t3779 (
    .I(seg_0_10_sp4_h_r_0_2238),
    .O(seg_0_12_sp4_v_b_24_2299)
  );
  CascadeMux t378 (
    .I(net_26993),
    .O(net_26993_cascademuxed)
  );
  Span4Mux_h4 t3780 (
    .I(seg_4_10_sp4_h_r_0_20174),
    .O(seg_0_10_sp4_h_r_0_2238)
  );
  Span4Mux_h4 t3781 (
    .I(seg_8_10_sp4_h_r_4_34873),
    .O(seg_4_10_sp4_h_r_0_20174)
  );
  LocalMux t3782 (
    .I(seg_8_10_sp4_h_r_8_34877),
    .O(seg_8_10_local_g0_0_34773)
  );
  LocalMux t3783 (
    .I(seg_9_15_sp4_r_v_b_11_38966),
    .O(seg_9_15_local_g2_3_39238)
  );
  Span4Mux_v4 t3784 (
    .I(seg_10_11_sp4_v_b_3_38466),
    .O(seg_9_15_sp4_r_v_b_11_38966)
  );
  LocalMux t3785 (
    .I(seg_10_15_sp4_v_b_11_38966),
    .O(seg_10_15_local_g1_3_43061)
  );
  Span4Mux_v4 t3786 (
    .I(seg_10_11_sp4_v_b_3_38466),
    .O(seg_10_15_sp4_v_b_11_38966)
  );
  LocalMux t3787 (
    .I(seg_9_15_sp4_r_v_b_22_39089),
    .O(seg_9_15_local_g3_6_39249)
  );
  Span4Mux_v3 t3788 (
    .I(seg_10_12_sp4_v_b_8_38596),
    .O(seg_9_15_sp4_r_v_b_22_39089)
  );
  LocalMux t3789 (
    .I(seg_10_15_sp4_v_b_22_39089),
    .O(seg_10_15_local_g0_6_43056)
  );
  Span4Mux_v3 t3790 (
    .I(seg_10_12_sp4_v_b_8_38596),
    .O(seg_10_15_sp4_v_b_22_39089)
  );
  LocalMux t3791 (
    .I(seg_10_7_sp4_v_b_41_38346),
    .O(seg_10_7_local_g3_1_42091)
  );
  LocalMux t3792 (
    .I(seg_9_12_sp4_r_v_b_22_38720),
    .O(seg_9_12_local_g3_6_38880)
  );
  LocalMux t3793 (
    .I(seg_10_11_lutff_0_out_38686),
    .O(seg_10_11_local_g0_0_42558)
  );
  LocalMux t3794 (
    .I(seg_11_12_neigh_op_bnl_1_38687),
    .O(seg_11_12_local_g2_1_46529)
  );
  LocalMux t3795 (
    .I(seg_10_11_lutff_3_out_38689),
    .O(seg_10_11_local_g1_3_42569)
  );
  LocalMux t3796 (
    .I(seg_11_11_neigh_op_lft_6_38692),
    .O(seg_11_11_local_g0_6_46395)
  );
  LocalMux t3797 (
    .I(seg_8_15_sp4_v_b_0_31295),
    .O(seg_8_15_local_g0_0_35388)
  );
  Span4Mux_v4 t3798 (
    .I(seg_8_11_sp4_h_r_0_34990),
    .O(seg_8_15_sp4_v_b_0_31295)
  );
  LocalMux t3799 (
    .I(seg_8_15_sp4_v_b_6_31301),
    .O(seg_8_15_local_g1_6_35402)
  );
  CascadeMux t38 (
    .I(net_8266),
    .O(net_8266_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t380 (
    .carryinitin(),
    .carryinitout(t379)
  );
  Span4Mux_v4 t3800 (
    .I(seg_8_11_sp4_h_r_6_34998),
    .O(seg_8_15_sp4_v_b_6_31301)
  );
  LocalMux t3801 (
    .I(seg_8_14_sp4_r_v_b_27_35250),
    .O(seg_8_14_local_g1_3_35276)
  );
  Span4Mux_v2 t3802 (
    .I(seg_9_12_sp4_h_r_9_38955),
    .O(seg_8_14_sp4_r_v_b_27_35250)
  );
  LocalMux t3803 (
    .I(seg_9_13_neigh_op_rgt_1_38933),
    .O(seg_9_13_local_g2_1_38990)
  );
  LocalMux t3804 (
    .I(seg_9_14_neigh_op_bnr_2_38934),
    .O(seg_9_14_local_g0_2_39098)
  );
  LocalMux t3805 (
    .I(seg_9_18_sp4_r_v_b_4_39330),
    .O(seg_9_18_local_g1_4_39600)
  );
  Span4Mux_v4 t3806 (
    .I(seg_10_14_sp4_h_r_10_43023),
    .O(seg_9_18_sp4_r_v_b_4_39330)
  );
  LocalMux t3807 (
    .I(seg_9_18_sp4_v_b_11_35504),
    .O(seg_9_18_local_g0_3_39591)
  );
  Span4Mux_v4 t3808 (
    .I(seg_9_14_sp4_h_r_5_39197),
    .O(seg_9_18_sp4_v_b_11_35504)
  );
  LocalMux t3809 (
    .I(seg_11_18_sp4_r_v_b_5_46991),
    .O(seg_11_18_local_g1_5_47263)
  );
  CascadeMux t381 (
    .I(net_27497),
    .O(net_27497_cascademuxed)
  );
  Span4Mux_v4 t3810 (
    .I(seg_12_14_sp4_h_l_37_35359),
    .O(seg_11_18_sp4_r_v_b_5_46991)
  );
  LocalMux t3811 (
    .I(seg_8_15_sp4_h_r_19_31659),
    .O(seg_8_15_local_g1_3_35399)
  );
  Span4Mux_h3 t3812 (
    .I(seg_11_15_sp4_v_b_6_42794),
    .O(seg_8_15_sp4_h_r_19_31659)
  );
  LocalMux t3813 (
    .I(seg_8_15_sp4_h_r_23_31653),
    .O(seg_8_15_local_g1_7_35403)
  );
  Span4Mux_h3 t3814 (
    .I(seg_11_15_sp4_v_b_10_42798),
    .O(seg_8_15_sp4_h_r_23_31653)
  );
  LocalMux t3815 (
    .I(seg_9_18_sp4_r_v_b_14_39450),
    .O(seg_9_18_local_g2_6_39610)
  );
  Span4Mux_v3 t3816 (
    .I(seg_10_15_sp4_v_b_3_38958),
    .O(seg_9_18_sp4_r_v_b_14_39450)
  );
  LocalMux t3817 (
    .I(seg_9_15_neigh_op_rgt_0_39178),
    .O(seg_9_15_local_g2_0_39235)
  );
  LocalMux t3818 (
    .I(seg_9_15_neigh_op_rgt_4_39182),
    .O(seg_9_15_local_g3_4_39247)
  );
  LocalMux t3819 (
    .I(seg_10_15_lutff_7_out_39185),
    .O(seg_10_15_local_g1_7_43065)
  );
  CascadeMux t382 (
    .I(net_27498),
    .O(net_27498_cascademuxed)
  );
  LocalMux t3820 (
    .I(seg_9_18_sp4_r_v_b_1_39325),
    .O(seg_9_18_local_g1_1_39597)
  );
  LocalMux t3821 (
    .I(seg_10_17_neigh_op_bot_0_39301),
    .O(seg_10_17_local_g0_0_43296)
  );
  LocalMux t3822 (
    .I(seg_9_17_neigh_op_bnr_1_39302),
    .O(seg_9_17_local_g1_1_39474)
  );
  LocalMux t3823 (
    .I(seg_9_17_neigh_op_bnr_3_39304),
    .O(seg_9_17_local_g1_3_39476)
  );
  LocalMux t3824 (
    .I(seg_10_17_neigh_op_bot_4_39305),
    .O(seg_10_17_local_g0_4_43300)
  );
  LocalMux t3825 (
    .I(seg_10_17_neigh_op_bot_5_39306),
    .O(seg_10_17_local_g0_5_43301)
  );
  LocalMux t3826 (
    .I(seg_9_18_neigh_op_bnr_0_39424),
    .O(seg_9_18_local_g1_0_39596)
  );
  LocalMux t3827 (
    .I(seg_9_18_neigh_op_bnr_1_39425),
    .O(seg_9_18_local_g0_1_39589)
  );
  LocalMux t3828 (
    .I(seg_9_18_neigh_op_bnr_2_39426),
    .O(seg_9_18_local_g0_2_39590)
  );
  LocalMux t3829 (
    .I(seg_9_18_neigh_op_bnr_4_39428),
    .O(seg_9_18_local_g0_4_39592)
  );
  LocalMux t3830 (
    .I(seg_9_18_neigh_op_bnr_6_39430),
    .O(seg_9_18_local_g1_6_39602)
  );
  LocalMux t3831 (
    .I(seg_9_18_neigh_op_bnr_7_39431),
    .O(seg_9_18_local_g0_7_39595)
  );
  LocalMux t3832 (
    .I(seg_10_18_lutff_1_out_39548),
    .O(seg_10_18_local_g1_1_43428)
  );
  LocalMux t3833 (
    .I(seg_10_18_lutff_2_out_39549),
    .O(seg_10_18_local_g2_2_43437)
  );
  LocalMux t3834 (
    .I(seg_10_18_lutff_3_out_39550),
    .O(seg_10_18_local_g2_3_43438)
  );
  LocalMux t3835 (
    .I(seg_10_18_lutff_5_out_39552),
    .O(seg_10_18_local_g3_5_43448)
  );
  LocalMux t3836 (
    .I(seg_10_18_lutff_6_out_39553),
    .O(seg_10_18_local_g2_6_43441)
  );
  LocalMux t3837 (
    .I(seg_10_18_lutff_7_out_39554),
    .O(seg_10_18_local_g0_7_43426)
  );
  LocalMux t3838 (
    .I(seg_14_18_sp4_h_r_8_58846),
    .O(seg_14_18_local_g0_0_58742)
  );
  Span4Mux_h0 t3839 (
    .I(seg_14_18_sp4_h_l_37_43513),
    .O(seg_14_18_sp4_h_r_8_58846)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t384 (
    .carryinitin(),
    .carryinitout(t383)
  );
  LocalMux t3840 (
    .I(seg_14_18_sp4_h_r_11_58839),
    .O(seg_14_18_local_g0_3_58745)
  );
  Span4Mux_h0 t3841 (
    .I(seg_14_18_sp4_h_l_45_43523),
    .O(seg_14_18_sp4_h_r_11_58839)
  );
  LocalMux t3842 (
    .I(seg_10_10_sp4_r_v_b_29_42422),
    .O(seg_10_10_local_g1_5_42448)
  );
  Span4Mux_v2 t3843 (
    .I(seg_11_12_sp4_v_t_39_42913),
    .O(seg_10_10_sp4_r_v_b_29_42422)
  );
  Span4Mux_v4 t3844 (
    .I(seg_11_16_sp4_v_t_39_43405),
    .O(seg_11_12_sp4_v_t_39_42913)
  );
  LocalMux t3845 (
    .I(seg_11_11_sp4_h_r_3_46488),
    .O(seg_11_11_local_g0_3_46392)
  );
  Span4Mux_h0 t3846 (
    .I(seg_11_11_sp4_v_t_38_42789),
    .O(seg_11_11_sp4_h_r_3_46488)
  );
  Span4Mux_v4 t3847 (
    .I(seg_11_15_sp4_v_t_38_43281),
    .O(seg_11_11_sp4_v_t_38_42789)
  );
  LocalMux t3848 (
    .I(seg_13_1_sp4_h_r_20_49059),
    .O(seg_13_1_local_g1_4_52793)
  );
  Span4Mux_h1 t3849 (
    .I(seg_12_1_sp4_v_b_9_45276),
    .O(seg_13_1_sp4_h_r_20_49059)
  );
  CascadeMux t385 (
    .I(net_27701),
    .O(net_27701_cascademuxed)
  );
  LocalMux t3850 (
    .I(seg_12_2_neigh_op_lft_2_41376),
    .O(seg_12_2_local_g1_2_49123)
  );
  LocalMux t3851 (
    .I(seg_12_3_neigh_op_bnl_4_41378),
    .O(seg_12_3_local_g2_4_49256)
  );
  LocalMux t3852 (
    .I(seg_11_3_neigh_op_bot_7_41381),
    .O(seg_11_3_local_g0_7_45412)
  );
  LocalMux t3853 (
    .I(seg_25_6_sp4_h_r_24_91207),
    .O(seg_25_6_local_g2_0_99386)
  );
  Span4Mux_h2 t3854 (
    .I(seg_23_6_sp4_v_b_6_87026),
    .O(seg_25_6_sp4_h_r_24_91207)
  );
  Span4Mux_v4 t3855 (
    .I(seg_23_2_sp4_h_l_43_75987),
    .O(seg_23_6_sp4_v_b_6_87026)
  );
  Span4Mux_h4 t3856 (
    .I(seg_19_2_sp4_h_l_43_60706),
    .O(seg_23_2_sp4_h_l_43_75987)
  );
  Span4Mux_h4 t3857 (
    .I(seg_15_2_sp4_h_l_47_45378),
    .O(seg_19_2_sp4_h_l_43_60706)
  );
  LocalMux t3858 (
    .I(seg_25_7_sp4_v_b_16_94983),
    .O(seg_25_7_local_g0_0_99520)
  );
  Span4Mux_v3 t3859 (
    .I(seg_25_4_sp4_v_b_2_90451),
    .O(seg_25_7_sp4_v_b_16_94983)
  );
  CascadeMux t386 (
    .I(net_27702),
    .O(net_27702_cascademuxed)
  );
  IoSpan4Mux t3860 (
    .I(seg_23_0_span4_vert_19_86748),
    .O(seg_25_4_sp4_v_b_2_90451)
  );
  Span4Mux_v2 t3861 (
    .I(seg_23_2_sp4_h_l_43_75987),
    .O(seg_23_0_span4_vert_19_86748)
  );
  LocalMux t3862 (
    .I(seg_13_4_sp4_v_b_33_49350),
    .O(seg_13_4_local_g2_1_53207)
  );
  Span4Mux_v2 t3863 (
    .I(seg_13_2_sp4_h_l_41_37720),
    .O(seg_13_4_sp4_v_b_33_49350)
  );
  LocalMux t3864 (
    .I(seg_13_4_sp4_v_b_27_49344),
    .O(seg_13_4_local_g3_3_53217)
  );
  Span4Mux_v2 t3865 (
    .I(seg_13_2_sp4_h_l_47_37716),
    .O(seg_13_4_sp4_v_b_27_49344)
  );
  LocalMux t3866 (
    .I(seg_11_4_neigh_op_bot_1_41534),
    .O(seg_11_4_local_g0_1_45529)
  );
  LocalMux t3867 (
    .I(seg_11_4_neigh_op_bot_2_41535),
    .O(seg_11_4_local_g1_2_45538)
  );
  LocalMux t3868 (
    .I(seg_11_4_neigh_op_bot_3_41536),
    .O(seg_11_4_local_g1_3_45539)
  );
  LocalMux t3869 (
    .I(seg_11_4_neigh_op_bot_4_41537),
    .O(seg_11_4_local_g0_4_45532)
  );
  CascadeMux t387 (
    .I(net_30116),
    .O(net_30116_cascademuxed)
  );
  LocalMux t3870 (
    .I(seg_11_4_neigh_op_bot_5_41538),
    .O(seg_11_4_local_g1_5_45541)
  );
  LocalMux t3871 (
    .I(seg_11_4_neigh_op_bot_6_41539),
    .O(seg_11_4_local_g1_6_45542)
  );
  LocalMux t3872 (
    .I(seg_11_4_neigh_op_bot_7_41540),
    .O(seg_11_4_local_g1_7_45543)
  );
  LocalMux t3873 (
    .I(seg_11_5_neigh_op_bot_3_41659),
    .O(seg_11_5_local_g1_3_45662)
  );
  LocalMux t3874 (
    .I(seg_12_3_neigh_op_tnl_5_41661),
    .O(seg_12_3_local_g2_5_49257)
  );
  LocalMux t3875 (
    .I(seg_13_4_sp12_h_r_10_34126),
    .O(seg_13_4_local_g1_2_53200)
  );
  LocalMux t3876 (
    .I(seg_13_3_sp4_v_b_23_49102),
    .O(seg_13_3_local_g0_7_53074)
  );
  Span4Mux_v1 t3877 (
    .I(seg_13_4_sp4_h_l_41_37966),
    .O(seg_13_3_sp4_v_b_23_49102)
  );
  LocalMux t3878 (
    .I(seg_13_4_sp4_h_r_32_45632),
    .O(seg_13_4_local_g2_0_53206)
  );
  LocalMux t3879 (
    .I(seg_12_2_sp4_v_b_29_45264),
    .O(seg_12_2_local_g2_5_49134)
  );
  CascadeMux t388 (
    .I(net_30269),
    .O(net_30269_cascademuxed)
  );
  LocalMux t3880 (
    .I(seg_11_2_sp4_v_b_38_41559),
    .O(seg_11_2_local_g2_6_45304)
  );
  LocalMux t3881 (
    .I(seg_11_2_sp4_v_b_26_41431),
    .O(seg_11_2_local_g2_2_45300)
  );
  LocalMux t3882 (
    .I(seg_10_6_neigh_op_bnr_2_41781),
    .O(seg_10_6_local_g1_2_41953)
  );
  LocalMux t3883 (
    .I(seg_12_4_neigh_op_tnl_3_41782),
    .O(seg_12_4_local_g2_3_49378)
  );
  LocalMux t3884 (
    .I(seg_11_5_lutff_6_out_41785),
    .O(seg_11_5_local_g1_6_45665)
  );
  LocalMux t3885 (
    .I(seg_13_5_sp4_h_r_34_45747),
    .O(seg_13_5_local_g2_2_53331)
  );
  LocalMux t3886 (
    .I(seg_15_5_sp4_h_r_1_61068),
    .O(seg_15_5_local_g1_1_60982)
  );
  Span4Mux_h0 t3887 (
    .I(seg_15_5_sp4_h_l_47_45747),
    .O(seg_15_5_sp4_h_r_1_61068)
  );
  LocalMux t3888 (
    .I(seg_13_6_sp4_v_b_39_49714),
    .O(seg_13_6_local_g3_7_53467)
  );
  Span4Mux_v1 t3889 (
    .I(seg_13_5_sp4_h_l_39_38087),
    .O(seg_13_6_sp4_v_b_39_49714)
  );
  CascadeMux t389 (
    .I(net_30281),
    .O(net_30281_cascademuxed)
  );
  LocalMux t3890 (
    .I(seg_14_4_sp4_r_v_b_23_56891),
    .O(seg_14_4_local_g3_7_57051)
  );
  Span4Mux_v1 t3891 (
    .I(seg_15_5_sp4_h_l_41_45751),
    .O(seg_14_4_sp4_r_v_b_23_56891)
  );
  LocalMux t3892 (
    .I(seg_14_5_sp4_h_r_41_45751),
    .O(seg_14_5_local_g3_1_57168)
  );
  LocalMux t3893 (
    .I(seg_15_5_sp4_h_r_7_61076),
    .O(seg_15_5_local_g1_7_60988)
  );
  Span4Mux_h0 t3894 (
    .I(seg_15_5_sp4_h_l_41_45751),
    .O(seg_15_5_sp4_h_r_7_61076)
  );
  LocalMux t3895 (
    .I(seg_12_7_sp4_v_b_19_45764),
    .O(seg_12_7_local_g1_3_49739)
  );
  LocalMux t3896 (
    .I(seg_12_8_sp4_v_b_6_45764),
    .O(seg_12_8_local_g0_6_49857)
  );
  LocalMux t3897 (
    .I(seg_11_2_sp4_v_b_37_41558),
    .O(seg_11_2_local_g3_5_45311)
  );
  LocalMux t3898 (
    .I(seg_11_3_sp4_v_b_38_41682),
    .O(seg_11_3_local_g2_6_45427)
  );
  LocalMux t3899 (
    .I(seg_11_2_sp4_v_b_39_41560),
    .O(seg_11_2_local_g3_7_45313)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t39 (
    .carryinitin(net_12615),
    .carryinitout(net_12659)
  );
  CascadeMux t390 (
    .I(net_30362),
    .O(net_30362_cascademuxed)
  );
  LocalMux t3900 (
    .I(seg_13_6_sp4_h_r_27_45873),
    .O(seg_13_6_local_g2_3_53455)
  );
  Span4Mux_h2 t3901 (
    .I(seg_11_6_sp4_v_b_9_41688),
    .O(seg_13_6_sp4_h_r_27_45873)
  );
  LocalMux t3902 (
    .I(seg_11_3_sp4_v_b_30_41564),
    .O(seg_11_3_local_g3_6_45435)
  );
  LocalMux t3903 (
    .I(seg_11_3_sp4_v_b_32_41566),
    .O(seg_11_3_local_g3_0_45429)
  );
  LocalMux t3904 (
    .I(seg_11_6_lutff_0_out_41902),
    .O(seg_11_6_local_g2_0_45790)
  );
  LocalMux t3905 (
    .I(seg_10_6_neigh_op_rgt_1_41903),
    .O(seg_10_6_local_g3_1_41968)
  );
  LocalMux t3906 (
    .I(seg_11_5_neigh_op_top_4_41906),
    .O(seg_11_5_local_g1_4_45663)
  );
  LocalMux t3907 (
    .I(seg_11_5_neigh_op_top_7_41909),
    .O(seg_11_5_local_g1_7_45666)
  );
  LocalMux t3908 (
    .I(seg_14_5_sp4_v_b_12_53173),
    .O(seg_14_5_local_g1_4_57155)
  );
  Span4Mux_v1 t3909 (
    .I(seg_14_6_sp4_h_l_42_42046),
    .O(seg_14_5_sp4_v_b_12_53173)
  );
  CascadeMux t391 (
    .I(net_30368),
    .O(net_30368_cascademuxed)
  );
  LocalMux t3910 (
    .I(seg_13_6_sp4_h_r_26_45872),
    .O(seg_13_6_local_g2_2_53454)
  );
  LocalMux t3911 (
    .I(seg_15_5_sp4_v_b_21_57012),
    .O(seg_15_5_local_g0_5_60978)
  );
  Span4Mux_v1 t3912 (
    .I(seg_15_6_sp4_h_l_39_45872),
    .O(seg_15_5_sp4_v_b_21_57012)
  );
  LocalMux t3913 (
    .I(seg_14_4_sp4_h_r_28_49459),
    .O(seg_14_4_local_g2_4_57040)
  );
  Span4Mux_h2 t3914 (
    .I(seg_12_4_sp4_v_t_46_45767),
    .O(seg_14_4_sp4_h_r_28_49459)
  );
  LocalMux t3915 (
    .I(seg_15_6_sp4_v_b_13_57127),
    .O(seg_15_6_local_g1_5_61109)
  );
  Span4Mux_v1 t3916 (
    .I(seg_15_7_sp4_h_l_37_45991),
    .O(seg_15_6_sp4_v_b_13_57127)
  );
  LocalMux t3917 (
    .I(seg_15_6_sp4_v_b_17_57131),
    .O(seg_15_6_local_g0_1_61097)
  );
  Span4Mux_v1 t3918 (
    .I(seg_15_7_sp4_h_l_47_45993),
    .O(seg_15_6_sp4_v_b_17_57131)
  );
  LocalMux t3919 (
    .I(seg_15_6_sp4_h_r_41_49705),
    .O(seg_15_6_local_g3_1_61121)
  );
  CascadeMux t392 (
    .I(net_30374),
    .O(net_30374_cascademuxed)
  );
  Span4Mux_h3 t3920 (
    .I(seg_12_6_sp4_v_t_41_46008),
    .O(seg_15_6_sp4_h_r_41_49705)
  );
  LocalMux t3921 (
    .I(seg_12_7_neigh_op_tnl_0_42148),
    .O(seg_12_7_local_g2_0_49744)
  );
  LocalMux t3922 (
    .I(seg_12_8_neigh_op_lft_0_42148),
    .O(seg_12_8_local_g1_0_49859)
  );
  LocalMux t3923 (
    .I(seg_11_8_lutff_1_out_42149),
    .O(seg_11_8_local_g0_1_46021)
  );
  LocalMux t3924 (
    .I(seg_12_8_neigh_op_lft_2_42150),
    .O(seg_12_8_local_g1_2_49861)
  );
  LocalMux t3925 (
    .I(seg_11_8_lutff_4_out_42152),
    .O(seg_11_8_local_g2_4_46040)
  );
  LocalMux t3926 (
    .I(seg_0_25_sp4_v_b_7_4668),
    .O(seg_0_25_local_g0_7_5328)
  );
  Span4Mux_v4 t3927 (
    .I(seg_0_21_sp4_h_r_1_4603),
    .O(seg_0_25_sp4_v_b_7_4668)
  );
  Span4Mux_h4 t3928 (
    .I(seg_4_21_sp4_v_b_1_17339),
    .O(seg_0_21_sp4_h_r_1_4603)
  );
  Sp12to4 t3929 (
    .I(seg_4_20_sp12_v_b_1_19926),
    .O(seg_4_21_sp4_v_b_1_17339)
  );
  CascadeMux t393 (
    .I(net_30380),
    .O(net_30380_cascademuxed)
  );
  Span12Mux_v12 t3930 (
    .I(seg_4_8_sp12_h_r_1_19925),
    .O(seg_4_20_sp12_v_b_1_19926)
  );
  LocalMux t3931 (
    .I(seg_0_25_sp4_r_v_b_12_5087),
    .O(seg_0_25_local_g2_4_5341)
  );
  Span4Mux_v3 t3932 (
    .I(seg_1_22_sp4_v_b_10_4207),
    .O(seg_0_25_sp4_r_v_b_12_5087)
  );
  Span4Mux_v4 t3933 (
    .I(seg_1_18_sp4_v_b_2_3349),
    .O(seg_1_22_sp4_v_b_10_4207)
  );
  Sp12to4 t3934 (
    .I(seg_1_17_sp12_v_b_7_7901),
    .O(seg_1_18_sp4_v_b_2_3349)
  );
  Span12Mux_v9 t3935 (
    .I(seg_1_8_sp12_h_r_0_7898),
    .O(seg_1_17_sp12_v_b_7_7901)
  );
  LocalMux t3936 (
    .I(seg_0_25_sp4_v_b_4_4667),
    .O(seg_0_25_local_g0_4_5325)
  );
  Span4Mux_v4 t3937 (
    .I(seg_0_21_sp4_v_b_1_3772),
    .O(seg_0_25_sp4_v_b_4_4667)
  );
  Sp12to4 t3938 (
    .I(seg_0_20_sp12_v_b_1_1787),
    .O(seg_0_21_sp4_v_b_1_3772)
  );
  Span12Mux_v12 t3939 (
    .I(seg_0_8_sp12_h_r_1_1764),
    .O(seg_0_20_sp12_v_b_1_1787)
  );
  CascadeMux t394 (
    .I(net_30386),
    .O(net_30386_cascademuxed)
  );
  LocalMux t3940 (
    .I(seg_0_25_sp12_h_r_2_5427),
    .O(seg_0_25_local_g0_2_5323)
  );
  Span12Mux_h11 t3941 (
    .I(seg_11_25_sp12_v_b_1_46727),
    .O(seg_0_25_sp12_h_r_2_5427)
  );
  Span12Mux_v12 t3942 (
    .I(seg_11_13_sp12_v_b_1_45215),
    .O(seg_11_25_sp12_v_b_1_46727)
  );
  LocalMux t3943 (
    .I(seg_13_6_sp4_r_v_b_27_53421),
    .O(seg_13_6_local_g0_3_53439)
  );
  Span4Mux_v2 t3944 (
    .I(seg_14_8_sp4_h_l_44_42294),
    .O(seg_13_6_sp4_r_v_b_27_53421)
  );
  LocalMux t3945 (
    .I(seg_0_12_sp4_v_b_1_1861),
    .O(seg_0_12_local_g0_1_2521)
  );
  Span4Mux_v4 t3946 (
    .I(seg_0_8_sp4_h_r_7_1846),
    .O(seg_0_12_sp4_v_b_1_1861)
  );
  Span4Mux_h4 t3947 (
    .I(seg_4_8_sp4_h_r_11_19931),
    .O(seg_0_8_sp4_h_r_7_1846)
  );
  Span4Mux_h4 t3948 (
    .I(seg_8_8_sp4_h_r_3_34626),
    .O(seg_4_8_sp4_h_r_11_19931)
  );
  LocalMux t3949 (
    .I(seg_0_12_sp4_v_b_4_1866),
    .O(seg_0_12_local_g0_4_2524)
  );
  CascadeMux t395 (
    .I(net_30392),
    .O(net_30392_cascademuxed)
  );
  Span4Mux_v4 t3950 (
    .I(seg_0_8_sp4_h_r_10_1803),
    .O(seg_0_12_sp4_v_b_4_1866)
  );
  Span4Mux_h4 t3951 (
    .I(seg_4_8_sp4_h_r_10_19930),
    .O(seg_0_8_sp4_h_r_10_1803)
  );
  Span4Mux_h4 t3952 (
    .I(seg_8_8_sp4_h_r_7_34630),
    .O(seg_4_8_sp4_h_r_10_19930)
  );
  LocalMux t3953 (
    .I(seg_0_12_sp4_v_b_7_1867),
    .O(seg_0_12_local_g1_7_2535)
  );
  Span4Mux_v4 t3954 (
    .I(seg_0_8_sp4_h_r_1_1802),
    .O(seg_0_12_sp4_v_b_7_1867)
  );
  Span4Mux_h4 t3955 (
    .I(seg_4_8_sp4_h_r_5_19935),
    .O(seg_0_8_sp4_h_r_1_1802)
  );
  Span4Mux_h4 t3956 (
    .I(seg_8_8_sp4_h_r_9_34632),
    .O(seg_4_8_sp4_h_r_5_19935)
  );
  LocalMux t3957 (
    .I(seg_0_12_sp4_v_b_8_1870),
    .O(seg_0_12_local_g0_0_2520)
  );
  Span4Mux_v4 t3958 (
    .I(seg_0_8_sp4_h_r_2_1813),
    .O(seg_0_12_sp4_v_b_8_1870)
  );
  Span4Mux_h4 t3959 (
    .I(seg_4_8_sp4_h_r_2_19932),
    .O(seg_0_8_sp4_h_r_2_1813)
  );
  CascadeMux t396 (
    .I(net_30398),
    .O(net_30398_cascademuxed)
  );
  Span4Mux_h4 t3960 (
    .I(seg_8_8_sp4_h_r_11_34624),
    .O(seg_4_8_sp4_h_r_2_19932)
  );
  LocalMux t3961 (
    .I(seg_13_5_sp4_h_r_17_49582),
    .O(seg_13_5_local_g1_1_53322)
  );
  Span4Mux_h1 t3962 (
    .I(seg_12_5_sp4_v_t_41_45885),
    .O(seg_13_5_sp4_h_r_17_49582)
  );
  LocalMux t3963 (
    .I(seg_15_5_sp4_h_r_41_49582),
    .O(seg_15_5_local_g3_1_60998)
  );
  Span4Mux_h3 t3964 (
    .I(seg_12_5_sp4_v_t_41_45885),
    .O(seg_15_5_sp4_h_r_41_49582)
  );
  LocalMux t3965 (
    .I(seg_14_5_sp4_h_r_32_49586),
    .O(seg_14_5_local_g2_0_57159)
  );
  Span4Mux_h2 t3966 (
    .I(seg_12_5_sp4_v_t_45_45889),
    .O(seg_14_5_sp4_h_r_32_49586)
  );
  LocalMux t3967 (
    .I(seg_15_5_sp4_h_r_36_49577),
    .O(seg_15_5_local_g2_4_60993)
  );
  Span4Mux_h3 t3968 (
    .I(seg_12_5_sp4_v_t_45_45889),
    .O(seg_15_5_sp4_h_r_36_49577)
  );
  LocalMux t3969 (
    .I(seg_13_6_sp4_h_r_15_49703),
    .O(seg_13_6_local_g1_7_53451)
  );
  CascadeMux t397 (
    .I(net_30485),
    .O(net_30485_cascademuxed)
  );
  Span4Mux_h1 t3970 (
    .I(seg_12_6_sp4_v_t_44_46011),
    .O(seg_13_6_sp4_h_r_15_49703)
  );
  LocalMux t3971 (
    .I(seg_14_4_sp4_h_r_44_45633),
    .O(seg_14_4_local_g3_4_57048)
  );
  Span4Mux_h3 t3972 (
    .I(seg_11_4_sp4_v_t_41_41931),
    .O(seg_14_4_sp4_h_r_44_45633)
  );
  LocalMux t3973 (
    .I(seg_11_9_lutff_1_out_42272),
    .O(seg_11_9_local_g0_1_46144)
  );
  LocalMux t3974 (
    .I(seg_11_10_neigh_op_bot_7_42278),
    .O(seg_11_10_local_g0_7_46273)
  );
  LocalMux t3975 (
    .I(seg_11_11_sp4_v_b_0_42296),
    .O(seg_11_11_local_g0_0_46389)
  );
  LocalMux t3976 (
    .I(seg_10_11_sp4_r_v_b_6_42302),
    .O(seg_10_11_local_g1_6_42572)
  );
  LocalMux t3977 (
    .I(seg_10_14_sp4_r_v_b_20_42795),
    .O(seg_10_14_local_g3_4_42955)
  );
  Span4Mux_v3 t3978 (
    .I(seg_11_11_sp4_v_b_6_42302),
    .O(seg_10_14_sp4_r_v_b_20_42795)
  );
  LocalMux t3979 (
    .I(seg_11_14_sp4_v_b_20_42795),
    .O(seg_11_14_local_g0_4_46762)
  );
  CascadeMux t398 (
    .I(net_30491),
    .O(net_30491_cascademuxed)
  );
  Span4Mux_v3 t3980 (
    .I(seg_11_11_sp4_v_b_6_42302),
    .O(seg_11_14_sp4_v_b_20_42795)
  );
  LocalMux t3981 (
    .I(seg_10_11_neigh_op_bnr_1_42395),
    .O(seg_10_11_local_g0_1_42559)
  );
  LocalMux t3982 (
    .I(seg_11_11_neigh_op_bot_4_42398),
    .O(seg_11_11_local_g1_4_46401)
  );
  LocalMux t3983 (
    .I(seg_10_11_neigh_op_bnr_7_42401),
    .O(seg_10_11_local_g0_7_42565)
  );
  LocalMux t3984 (
    .I(seg_11_11_lutff_1_out_42518),
    .O(seg_11_11_local_g3_1_46414)
  );
  LocalMux t3985 (
    .I(seg_11_11_lutff_4_out_42521),
    .O(seg_11_11_local_g2_4_46409)
  );
  LocalMux t3986 (
    .I(seg_11_11_lutff_5_out_42522),
    .O(seg_11_11_local_g2_5_46410)
  );
  LocalMux t3987 (
    .I(seg_11_11_lutff_6_out_42523),
    .O(seg_11_11_local_g1_6_46403)
  );
  LocalMux t3988 (
    .I(seg_0_25_sp4_v_b_14_4891),
    .O(seg_0_25_local_g0_6_5327)
  );
  Span4Mux_v3 t3989 (
    .I(seg_0_22_sp4_v_b_3_3983),
    .O(seg_0_25_sp4_v_b_14_4891)
  );
  CascadeMux t399 (
    .I(net_30497),
    .O(net_30497_cascademuxed)
  );
  Sp12to4 t3990 (
    .I(seg_0_21_sp12_v_b_5_2430),
    .O(seg_0_22_sp4_v_b_3_3983)
  );
  Span12Mux_v10 t3991 (
    .I(seg_0_11_sp12_h_r_1_2407),
    .O(seg_0_21_sp12_v_b_5_2430)
  );
  LocalMux t3992 (
    .I(seg_0_25_sp4_r_v_b_15_5090),
    .O(seg_0_25_local_g2_7_5344)
  );
  Span4Mux_v3 t3993 (
    .I(seg_1_22_sp4_h_r_2_9964),
    .O(seg_0_25_sp4_r_v_b_15_5090)
  );
  Sp12to4 t3994 (
    .I(seg_2_22_sp12_h_r_6_4803),
    .O(seg_1_22_sp4_h_r_2_9964)
  );
  Span12Mux_h9 t3995 (
    .I(seg_11_22_sp12_v_b_1_46358),
    .O(seg_2_22_sp12_h_r_6_4803)
  );
  LocalMux t3996 (
    .I(seg_0_25_sp12_h_r_3_5432),
    .O(seg_0_25_local_g1_3_5332)
  );
  Span12Mux_h11 t3997 (
    .I(seg_11_25_sp12_v_b_0_46728),
    .O(seg_0_25_sp12_h_r_3_5432)
  );
  Span12Mux_v12 t3998 (
    .I(seg_11_13_sp12_v_b_0_45216),
    .O(seg_11_25_sp12_v_b_0_46728)
  );
  LocalMux t3999 (
    .I(seg_13_18_sp4_r_v_b_19_54779),
    .O(seg_13_18_local_g3_3_54939)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t4 (
    .carryinitin(),
    .carryinitout(t3)
  );
  CascadeMux t40 (
    .I(net_8560),
    .O(net_8560_cascademuxed)
  );
  CascadeMux t400 (
    .I(net_30521),
    .O(net_30521_cascademuxed)
  );
  Span4Mux_v3 t4000 (
    .I(seg_14_15_sp4_v_b_10_54291),
    .O(seg_13_18_sp4_r_v_b_19_54779)
  );
  Span4Mux_v4 t4001 (
    .I(seg_14_11_sp4_h_l_40_42659),
    .O(seg_14_15_sp4_v_b_10_54291)
  );
  LocalMux t4002 (
    .I(seg_0_12_sp4_h_r_10_2654),
    .O(seg_0_12_local_g0_2_2522)
  );
  Span4Mux_h4 t4003 (
    .I(seg_4_12_sp4_h_r_2_20424),
    .O(seg_0_12_sp4_h_r_10_2654)
  );
  Span4Mux_h4 t4004 (
    .I(seg_8_12_sp4_h_r_2_35117),
    .O(seg_4_12_sp4_h_r_2_20424)
  );
  Span4Mux_h4 t4005 (
    .I(seg_12_12_sp4_v_b_2_46252),
    .O(seg_8_12_sp4_h_r_2_35117)
  );
  LocalMux t4006 (
    .I(seg_0_12_sp4_h_r_11_2655),
    .O(seg_0_12_local_g1_3_2531)
  );
  Span4Mux_h4 t4007 (
    .I(seg_4_12_sp4_h_r_8_20430),
    .O(seg_0_12_sp4_h_r_11_2655)
  );
  Span4Mux_h4 t4008 (
    .I(seg_8_12_sp4_h_r_8_35123),
    .O(seg_4_12_sp4_h_r_8_20430)
  );
  Span4Mux_h4 t4009 (
    .I(seg_12_12_sp4_v_b_8_46258),
    .O(seg_8_12_sp4_h_r_8_35123)
  );
  CascadeMux t401 (
    .I(net_30608),
    .O(net_30608_cascademuxed)
  );
  LocalMux t4010 (
    .I(seg_0_12_sp4_h_r_2_2664),
    .O(seg_0_12_local_g1_2_2530)
  );
  Span4Mux_h4 t4011 (
    .I(seg_4_12_sp4_h_r_6_20428),
    .O(seg_0_12_sp4_h_r_2_2664)
  );
  Span4Mux_h4 t4012 (
    .I(seg_8_12_sp4_h_r_10_35115),
    .O(seg_4_12_sp4_h_r_6_20428)
  );
  Span4Mux_h4 t4013 (
    .I(seg_12_12_sp4_v_b_10_46260),
    .O(seg_8_12_sp4_h_r_10_35115)
  );
  LocalMux t4014 (
    .I(seg_11_12_lutff_2_out_42642),
    .O(seg_11_12_local_g1_2_46522)
  );
  LocalMux t4015 (
    .I(seg_11_16_sp12_v_b_2_45743),
    .O(seg_11_16_local_g3_2_47030)
  );
  LocalMux t4016 (
    .I(seg_11_16_sp4_v_b_8_42919),
    .O(seg_11_16_local_g1_0_47012)
  );
  Span4Mux_v4 t4017 (
    .I(seg_11_12_sp4_h_r_2_46610),
    .O(seg_11_16_sp4_v_b_8_42919)
  );
  LocalMux t4018 (
    .I(seg_13_8_sp4_h_r_12_49946),
    .O(seg_13_8_local_g0_4_53686)
  );
  Span4Mux_h1 t4019 (
    .I(seg_12_8_sp4_v_t_36_46249),
    .O(seg_13_8_sp4_h_r_12_49946)
  );
  CascadeMux t402 (
    .I(net_30614),
    .O(net_30614_cascademuxed)
  );
  LocalMux t4020 (
    .I(seg_11_18_sp4_v_b_16_43283),
    .O(seg_11_18_local_g0_0_47250)
  );
  Span4Mux_v3 t4021 (
    .I(seg_11_15_sp4_v_b_5_42791),
    .O(seg_11_18_sp4_v_b_16_43283)
  );
  LocalMux t4022 (
    .I(seg_11_13_lutff_4_out_42767),
    .O(seg_11_13_local_g2_4_46655)
  );
  LocalMux t4023 (
    .I(seg_11_18_sp4_v_b_9_43164),
    .O(seg_11_18_local_g0_1_47251)
  );
  Span4Mux_v4 t4024 (
    .I(seg_11_14_sp4_v_b_9_42672),
    .O(seg_11_18_sp4_v_b_9_43164)
  );
  LocalMux t4025 (
    .I(seg_11_18_sp12_v_b_6_46235),
    .O(seg_11_18_local_g3_6_47280)
  );
  LocalMux t4026 (
    .I(seg_11_18_sp12_v_b_0_45867),
    .O(seg_11_18_local_g2_0_47266)
  );
  LocalMux t4027 (
    .I(seg_11_18_sp4_v_b_6_43163),
    .O(seg_11_18_local_g0_6_47256)
  );
  Span4Mux_v4 t4028 (
    .I(seg_11_14_sp4_h_r_0_46852),
    .O(seg_11_18_sp4_v_b_6_43163)
  );
  LocalMux t4029 (
    .I(seg_8_15_sp4_v_b_42_31669),
    .O(seg_8_15_local_g3_2_35414)
  );
  CascadeMux t403 (
    .I(net_30632),
    .O(net_30632_cascademuxed)
  );
  Span4Mux_v1 t4030 (
    .I(seg_8_14_sp4_h_r_7_35368),
    .O(seg_8_15_sp4_v_b_42_31669)
  );
  LocalMux t4031 (
    .I(seg_8_15_sp4_h_r_1_35483),
    .O(seg_8_15_local_g1_1_35397)
  );
  Span4Mux_h4 t4032 (
    .I(seg_12_15_sp4_v_b_8_46627),
    .O(seg_8_15_sp4_h_r_1_35483)
  );
  LocalMux t4033 (
    .I(seg_11_15_lutff_0_out_43009),
    .O(seg_11_15_local_g2_0_46897)
  );
  LocalMux t4034 (
    .I(seg_11_15_lutff_6_out_43015),
    .O(seg_11_15_local_g0_6_46887)
  );
  LocalMux t4035 (
    .I(seg_8_15_sp4_h_r_11_35485),
    .O(seg_8_15_local_g0_3_35391)
  );
  LocalMux t4036 (
    .I(seg_11_17_sp4_v_b_0_43034),
    .O(seg_11_17_local_g1_0_47135)
  );
  LocalMux t4037 (
    .I(seg_11_17_sp4_v_b_10_43044),
    .O(seg_11_17_local_g0_2_47129)
  );
  LocalMux t4038 (
    .I(seg_13_18_sp4_h_r_25_47345),
    .O(seg_13_18_local_g2_1_54929)
  );
  Span4Mux_h2 t4039 (
    .I(seg_11_18_sp4_v_b_1_43156),
    .O(seg_13_18_sp4_h_r_25_47345)
  );
  LocalMux t4040 (
    .I(seg_11_16_lutff_3_out_43135),
    .O(seg_11_16_local_g2_3_47023)
  );
  LocalMux t4041 (
    .I(seg_11_16_lutff_4_out_43136),
    .O(seg_11_16_local_g0_4_47008)
  );
  LocalMux t4042 (
    .I(seg_10_18_sp4_v_b_31_39577),
    .O(seg_10_18_local_g3_7_43450)
  );
  Span4Mux_v2 t4043 (
    .I(seg_10_16_sp4_h_r_7_43276),
    .O(seg_10_18_sp4_v_b_31_39577)
  );
  LocalMux t4044 (
    .I(seg_10_18_sp4_r_v_b_8_43165),
    .O(seg_10_18_local_g2_0_43435)
  );
  LocalMux t4045 (
    .I(seg_11_17_lutff_0_out_43255),
    .O(seg_11_17_local_g2_0_47143)
  );
  LocalMux t4046 (
    .I(seg_11_17_lutff_2_out_43257),
    .O(seg_11_17_local_g1_2_47137)
  );
  LocalMux t4047 (
    .I(seg_10_17_neigh_op_rgt_3_43258),
    .O(seg_10_17_local_g2_3_43315)
  );
  LocalMux t4048 (
    .I(seg_10_17_neigh_op_rgt_4_43259),
    .O(seg_10_17_local_g2_4_43316)
  );
  LocalMux t4049 (
    .I(seg_11_18_neigh_op_bot_5_43260),
    .O(seg_11_18_local_g0_5_47255)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t405 (
    .carryinitin(),
    .carryinitout(t404)
  );
  LocalMux t4050 (
    .I(seg_11_18_neigh_op_bot_6_43261),
    .O(seg_11_18_local_g1_6_47264)
  );
  LocalMux t4051 (
    .I(seg_10_17_neigh_op_rgt_7_43262),
    .O(seg_10_17_local_g2_7_43319)
  );
  LocalMux t4052 (
    .I(seg_10_18_neigh_op_rgt_1_43379),
    .O(seg_10_18_local_g3_1_43444)
  );
  LocalMux t4053 (
    .I(seg_11_12_sp4_r_v_b_47_46629),
    .O(seg_11_12_local_g3_7_46543)
  );
  Span4Mux_v3 t4054 (
    .I(seg_12_15_sp4_v_t_39_47113),
    .O(seg_11_12_sp4_r_v_b_47_46629)
  );
  LocalMux t4055 (
    .I(seg_11_16_sp4_r_v_b_45_47119),
    .O(seg_11_16_local_g3_5_47033)
  );
  LocalMux t4056 (
    .I(seg_12_14_sp4_v_b_30_46748),
    .O(seg_12_14_local_g3_6_50619)
  );
  Span4Mux_v2 t4057 (
    .I(seg_12_16_sp4_v_t_38_47235),
    .O(seg_12_14_sp4_v_b_30_46748)
  );
  LocalMux t4058 (
    .I(seg_10_19_neigh_op_rgt_1_43502),
    .O(seg_10_19_local_g2_1_43559)
  );
  LocalMux t4059 (
    .I(seg_11_2_neigh_op_bnr_1_45078),
    .O(seg_11_2_local_g0_1_45283)
  );
  CascadeMux t406 (
    .I(net_30743),
    .O(net_30743_cascademuxed)
  );
  LocalMux t4060 (
    .I(seg_12_1_lutff_1_out_45078),
    .O(seg_12_1_local_g1_1_48959)
  );
  LocalMux t4061 (
    .I(seg_12_1_lutff_2_out_45079),
    .O(seg_12_1_local_g0_2_48952)
  );
  LocalMux t4062 (
    .I(seg_12_2_neigh_op_bot_2_45079),
    .O(seg_12_2_local_g0_2_49115)
  );
  LocalMux t4063 (
    .I(seg_13_2_neigh_op_bnl_2_45079),
    .O(seg_13_2_local_g3_2_52970)
  );
  LocalMux t4064 (
    .I(seg_12_1_lutff_3_out_45080),
    .O(seg_12_1_local_g3_3_48977)
  );
  LocalMux t4065 (
    .I(seg_12_2_neigh_op_bot_3_45080),
    .O(seg_12_2_local_g1_3_49124)
  );
  LocalMux t4066 (
    .I(seg_13_2_neigh_op_bnl_3_45080),
    .O(seg_13_2_local_g3_3_52971)
  );
  LocalMux t4067 (
    .I(seg_12_1_lutff_4_out_45081),
    .O(seg_12_1_local_g0_4_48954)
  );
  LocalMux t4068 (
    .I(seg_14_2_sp4_h_r_19_53046),
    .O(seg_14_2_local_g1_3_56785)
  );
  Span4Mux_h1 t4069 (
    .I(seg_13_2_sp4_v_b_6_49071),
    .O(seg_14_2_sp4_h_r_19_53046)
  );
  CascadeMux t407 (
    .I(net_30755),
    .O(net_30755_cascademuxed)
  );
  LocalMux t4070 (
    .I(seg_14_2_sp4_h_r_21_53048),
    .O(seg_14_2_local_g0_5_56779)
  );
  Span4Mux_h1 t4071 (
    .I(seg_13_2_sp4_v_b_8_49074),
    .O(seg_14_2_sp4_h_r_21_53048)
  );
  LocalMux t4072 (
    .I(seg_14_2_sp4_h_r_17_53044),
    .O(seg_14_2_local_g1_1_56783)
  );
  Span4Mux_h1 t4073 (
    .I(seg_13_2_sp4_v_b_10_49076),
    .O(seg_14_2_sp4_h_r_17_53044)
  );
  LocalMux t4074 (
    .I(seg_14_3_sp4_h_r_18_53170),
    .O(seg_14_3_local_g1_2_56907)
  );
  Span4Mux_h1 t4075 (
    .I(seg_13_3_sp4_v_b_1_49078),
    .O(seg_14_3_sp4_h_r_18_53170)
  );
  LocalMux t4076 (
    .I(seg_13_3_sp4_v_b_11_49089),
    .O(seg_13_3_local_g0_3_53070)
  );
  LocalMux t4077 (
    .I(seg_13_4_sp4_v_b_0_49091),
    .O(seg_13_4_local_g1_0_53198)
  );
  LocalMux t4078 (
    .I(seg_13_4_sp4_v_b_2_49093),
    .O(seg_13_4_local_g0_2_53192)
  );
  LocalMux t4079 (
    .I(seg_12_4_sp4_r_v_b_4_49096),
    .O(seg_12_4_local_g1_4_49371)
  );
  CascadeMux t408 (
    .I(net_30896),
    .O(net_30896_cascademuxed)
  );
  LocalMux t4080 (
    .I(seg_13_3_sp4_v_b_17_49096),
    .O(seg_13_3_local_g0_1_53068)
  );
  LocalMux t4081 (
    .I(seg_13_4_sp4_v_b_4_49096),
    .O(seg_13_4_local_g0_4_53194)
  );
  LocalMux t4082 (
    .I(seg_12_3_sp4_v_b_10_45257),
    .O(seg_12_3_local_g0_2_49238)
  );
  LocalMux t4083 (
    .I(seg_12_3_neigh_op_bot_0_45205),
    .O(seg_12_3_local_g0_0_49236)
  );
  LocalMux t4084 (
    .I(seg_12_3_neigh_op_bot_2_45207),
    .O(seg_12_3_local_g1_2_49246)
  );
  LocalMux t4085 (
    .I(seg_11_2_neigh_op_rgt_3_45208),
    .O(seg_11_2_local_g2_3_45301)
  );
  LocalMux t4086 (
    .I(seg_12_2_lutff_6_out_45211),
    .O(seg_12_2_local_g0_6_49119)
  );
  LocalMux t4087 (
    .I(seg_15_2_sp4_h_r_39_49211),
    .O(seg_15_2_local_g2_7_60627)
  );
  LocalMux t4088 (
    .I(seg_15_4_sp4_r_v_b_26_60836),
    .O(seg_15_4_local_g1_2_60860)
  );
  Span4Mux_v2 t4089 (
    .I(seg_16_2_sp4_h_l_39_49211),
    .O(seg_15_4_sp4_r_v_b_26_60836)
  );
  CascadeMux t409 (
    .I(net_30983),
    .O(net_30983_cascademuxed)
  );
  LocalMux t4090 (
    .I(seg_16_2_sp4_h_r_5_64536),
    .O(seg_16_2_local_g0_5_64440)
  );
  Span4Mux_h0 t4091 (
    .I(seg_16_2_sp4_h_l_39_49211),
    .O(seg_16_2_sp4_h_r_5_64536)
  );
  LocalMux t4092 (
    .I(seg_9_2_sp4_h_r_3_37719),
    .O(seg_9_2_local_g1_3_37631)
  );
  LocalMux t4093 (
    .I(seg_14_4_sp4_h_r_12_53285),
    .O(seg_14_4_local_g1_4_57032)
  );
  Span4Mux_h1 t4094 (
    .I(seg_13_4_sp4_v_b_1_49090),
    .O(seg_14_4_sp4_h_r_12_53285)
  );
  LocalMux t4095 (
    .I(seg_14_5_sp4_h_r_17_53413),
    .O(seg_14_5_local_g1_1_57152)
  );
  Span4Mux_h1 t4096 (
    .I(seg_13_5_sp4_v_b_4_49224),
    .O(seg_14_5_sp4_h_r_17_53413)
  );
  LocalMux t4097 (
    .I(seg_15_5_sp4_h_r_28_53413),
    .O(seg_15_5_local_g3_4_61001)
  );
  Span4Mux_h2 t4098 (
    .I(seg_13_5_sp4_v_b_4_49224),
    .O(seg_15_5_sp4_h_r_28_53413)
  );
  LocalMux t4099 (
    .I(seg_8_7_sp4_v_b_5_30314),
    .O(seg_8_7_local_g0_5_34409)
  );
  CascadeMux t410 (
    .I(net_31001),
    .O(net_31001_cascademuxed)
  );
  Span4Mux_v4 t4100 (
    .I(seg_8_3_sp4_h_r_11_34009),
    .O(seg_8_7_sp4_v_b_5_30314)
  );
  Span4Mux_h4 t4101 (
    .I(seg_12_3_sp4_v_b_11_45258),
    .O(seg_8_3_sp4_h_r_11_34009)
  );
  LocalMux t4102 (
    .I(seg_9_3_sp4_h_r_22_34009),
    .O(seg_9_3_local_g0_6_37749)
  );
  Span4Mux_h3 t4103 (
    .I(seg_12_3_sp4_v_b_11_45258),
    .O(seg_9_3_sp4_h_r_22_34009)
  );
  LocalMux t4104 (
    .I(seg_9_4_sp4_h_r_14_34134),
    .O(seg_9_4_local_g0_6_37872)
  );
  Span4Mux_h3 t4105 (
    .I(seg_12_4_sp4_v_b_10_45271),
    .O(seg_9_4_sp4_h_r_14_34134)
  );
  LocalMux t4106 (
    .I(seg_10_4_sp4_h_r_27_34134),
    .O(seg_10_4_local_g3_3_41724)
  );
  Span4Mux_h2 t4107 (
    .I(seg_12_4_sp4_v_b_10_45271),
    .O(seg_10_4_sp4_h_r_27_34134)
  );
  LocalMux t4108 (
    .I(seg_12_5_sp4_v_b_3_45390),
    .O(seg_12_5_local_g1_3_49493)
  );
  LocalMux t4109 (
    .I(seg_12_5_sp4_v_b_5_45392),
    .O(seg_12_5_local_g1_5_49495)
  );
  CascadeMux t411 (
    .I(net_31100),
    .O(net_31100_cascademuxed)
  );
  LocalMux t4110 (
    .I(seg_12_8_sp4_v_b_12_45880),
    .O(seg_12_8_local_g0_4_49855)
  );
  Span4Mux_v3 t4111 (
    .I(seg_12_5_sp4_v_b_5_45392),
    .O(seg_12_8_sp4_v_b_12_45880)
  );
  LocalMux t4112 (
    .I(seg_12_3_lutff_4_out_45368),
    .O(seg_12_3_local_g0_4_49240)
  );
  LocalMux t4113 (
    .I(seg_12_4_neigh_op_bot_4_45368),
    .O(seg_12_4_local_g0_4_49363)
  );
  LocalMux t4114 (
    .I(seg_12_3_lutff_5_out_45369),
    .O(seg_12_3_local_g0_5_49241)
  );
  LocalMux t4115 (
    .I(seg_12_4_neigh_op_bot_6_45370),
    .O(seg_12_4_local_g0_6_49365)
  );
  LocalMux t4116 (
    .I(seg_0_25_sp4_v_b_13_4890),
    .O(seg_0_25_local_g0_5_5326)
  );
  Span4Mux_v3 t4117 (
    .I(seg_0_22_sp4_h_r_0_4829),
    .O(seg_0_25_sp4_v_b_13_4890)
  );
  Sp12to4 t4118 (
    .I(seg_1_22_sp12_h_r_2_4792),
    .O(seg_0_22_sp4_h_r_0_4829)
  );
  Span12Mux_h11 t4119 (
    .I(seg_12_22_sp12_v_b_1_50189),
    .O(seg_1_22_sp12_h_r_2_4792)
  );
  Span12Mux_v12 t4120 (
    .I(seg_12_10_sp12_v_b_1_48926),
    .O(seg_12_22_sp12_v_b_1_50189)
  );
  LocalMux t4121 (
    .I(seg_7_7_sp4_h_r_22_27322),
    .O(seg_7_7_local_g0_6_30579)
  );
  Span4Mux_h3 t4122 (
    .I(seg_10_7_sp4_v_b_6_37979),
    .O(seg_7_7_sp4_h_r_22_27322)
  );
  Span4Mux_v4 t4123 (
    .I(seg_10_3_sp4_h_r_0_41668),
    .O(seg_10_7_sp4_v_b_6_37979)
  );
  LocalMux t4124 (
    .I(seg_10_7_sp4_v_b_6_37979),
    .O(seg_10_7_local_g0_6_42072)
  );
  LocalMux t4125 (
    .I(seg_10_10_sp4_v_b_20_38472),
    .O(seg_10_10_local_g0_4_42439)
  );
  Span4Mux_v3 t4126 (
    .I(seg_10_7_sp4_v_b_6_37979),
    .O(seg_10_10_sp4_v_b_20_38472)
  );
  LocalMux t4127 (
    .I(seg_17_2_sp4_r_v_b_18_68238),
    .O(seg_17_2_local_g3_2_68292)
  );
  Span4Mux_v1 t4128 (
    .I(seg_18_3_sp4_h_l_42_57000),
    .O(seg_17_2_sp4_r_v_b_18_68238)
  );
  Span4Mux_h4 t4129 (
    .I(seg_14_3_sp4_h_l_41_41674),
    .O(seg_18_3_sp4_h_l_42_57000)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t413 (
    .carryinitin(),
    .carryinitout(t412)
  );
  LocalMux t4130 (
    .I(seg_4_6_sp4_r_v_b_16_19452),
    .O(seg_4_6_local_g3_0_19612)
  );
  Span4Mux_v3 t4131 (
    .I(seg_5_3_sp4_h_r_5_23151),
    .O(seg_4_6_sp4_r_v_b_16_19452)
  );
  Span4Mux_h4 t4132 (
    .I(seg_9_3_sp4_h_r_5_37844),
    .O(seg_5_3_sp4_h_r_5_23151)
  );
  LocalMux t4133 (
    .I(seg_5_4_sp4_v_b_40_19452),
    .O(seg_5_4_local_g3_0_23197)
  );
  Span4Mux_v1 t4134 (
    .I(seg_5_3_sp4_h_r_5_23151),
    .O(seg_5_4_sp4_v_b_40_19452)
  );
  LocalMux t4135 (
    .I(seg_9_7_sp4_v_b_5_34145),
    .O(seg_9_7_local_g0_5_38240)
  );
  Span4Mux_v4 t4136 (
    .I(seg_9_3_sp4_h_r_5_37844),
    .O(seg_9_7_sp4_v_b_5_34145)
  );
  LocalMux t4137 (
    .I(seg_9_10_sp4_v_b_12_34633),
    .O(seg_9_10_local_g1_4_38616)
  );
  Span4Mux_v3 t4138 (
    .I(seg_9_7_sp4_v_b_5_34145),
    .O(seg_9_10_sp4_v_b_12_34633)
  );
  LocalMux t4139 (
    .I(seg_11_11_sp4_r_v_b_5_46130),
    .O(seg_11_11_local_g1_5_46402)
  );
  Span4Mux_v4 t4140 (
    .I(seg_12_7_sp4_v_b_2_45637),
    .O(seg_11_11_sp4_r_v_b_5_46130)
  );
  Span4Mux_v4 t4141 (
    .I(seg_12_3_sp4_h_r_8_49340),
    .O(seg_12_7_sp4_v_b_2_45637)
  );
  LocalMux t4142 (
    .I(seg_5_8_sp4_v_b_15_19697),
    .O(seg_5_8_local_g0_7_23672)
  );
  Span4Mux_v3 t4143 (
    .I(seg_5_5_sp4_h_r_2_23394),
    .O(seg_5_8_sp4_v_b_15_19697)
  );
  Span4Mux_h4 t4144 (
    .I(seg_9_5_sp4_h_r_6_38091),
    .O(seg_5_5_sp4_h_r_2_23394)
  );
  Span4Mux_h4 t4145 (
    .I(seg_13_5_sp4_v_b_1_49219),
    .O(seg_9_5_sp4_h_r_6_38091)
  );
  LocalMux t4146 (
    .I(seg_12_5_sp4_r_v_b_21_49351),
    .O(seg_12_5_local_g3_5_49511)
  );
  LocalMux t4147 (
    .I(seg_10_4_sp4_h_r_30_34137),
    .O(seg_10_4_local_g2_6_41719)
  );
  Span4Mux_h2 t4148 (
    .I(seg_12_4_sp4_v_b_1_45259),
    .O(seg_10_4_sp4_h_r_30_34137)
  );
  LocalMux t4149 (
    .I(seg_15_4_sp4_h_r_42_49462),
    .O(seg_15_4_local_g3_2_60876)
  );
  Span4Mux_h3 t4150 (
    .I(seg_12_4_sp4_v_b_1_45259),
    .O(seg_15_4_sp4_h_r_42_49462)
  );
  LocalMux t4151 (
    .I(seg_4_5_sp4_h_r_1_19560),
    .O(seg_4_5_local_g1_1_19474)
  );
  Span4Mux_h4 t4152 (
    .I(seg_8_5_sp4_h_r_5_34259),
    .O(seg_4_5_sp4_h_r_1_19560)
  );
  Span4Mux_h4 t4153 (
    .I(seg_12_5_sp4_v_b_0_45389),
    .O(seg_8_5_sp4_h_r_5_34259)
  );
  LocalMux t4154 (
    .I(seg_7_4_sp4_r_v_b_23_30075),
    .O(seg_7_4_local_g3_7_30235)
  );
  Span4Mux_v1 t4155 (
    .I(seg_8_5_sp4_h_r_5_34259),
    .O(seg_7_4_sp4_r_v_b_23_30075)
  );
  LocalMux t4156 (
    .I(seg_8_5_sp4_h_r_5_34259),
    .O(seg_8_5_local_g1_5_34171)
  );
  LocalMux t4157 (
    .I(seg_9_5_sp4_h_r_16_34259),
    .O(seg_9_5_local_g0_0_37989)
  );
  Span4Mux_h3 t4158 (
    .I(seg_12_5_sp4_v_b_0_45389),
    .O(seg_9_5_sp4_h_r_16_34259)
  );
  LocalMux t4159 (
    .I(seg_11_8_sp4_r_v_b_14_45882),
    .O(seg_11_8_local_g2_6_46042)
  );
  Span4Mux_v3 t4160 (
    .I(seg_12_5_sp4_v_b_0_45389),
    .O(seg_11_8_sp4_r_v_b_14_45882)
  );
  LocalMux t4161 (
    .I(seg_12_16_sp4_v_b_20_46872),
    .O(seg_12_16_local_g0_4_50839)
  );
  Span4Mux_v3 t4162 (
    .I(seg_12_13_sp4_v_b_6_46379),
    .O(seg_12_16_sp4_v_b_20_46872)
  );
  Span4Mux_v4 t4163 (
    .I(seg_12_9_sp4_v_b_3_45882),
    .O(seg_12_13_sp4_v_b_6_46379)
  );
  Span4Mux_v4 t4164 (
    .I(seg_12_5_sp4_v_b_0_45389),
    .O(seg_12_9_sp4_v_b_3_45882)
  );
  LocalMux t4165 (
    .I(seg_0_12_sp4_v_b_19_2095),
    .O(seg_0_12_local_g0_3_2523)
  );
  Span4Mux_v3 t4166 (
    .I(seg_0_9_sp4_h_r_6_2072),
    .O(seg_0_12_sp4_v_b_19_2095)
  );
  Span4Mux_h4 t4167 (
    .I(seg_4_9_sp4_h_r_6_20059),
    .O(seg_0_9_sp4_h_r_6_2072)
  );
  Span4Mux_h4 t4168 (
    .I(seg_8_9_sp4_h_r_6_34752),
    .O(seg_4_9_sp4_h_r_6_20059)
  );
  Span4Mux_h4 t4169 (
    .I(seg_12_9_sp4_v_b_6_45887),
    .O(seg_8_9_sp4_h_r_6_34752)
  );
  Span4Mux_v4 t4170 (
    .I(seg_12_5_sp4_v_b_6_45395),
    .O(seg_12_9_sp4_v_b_6_45887)
  );
  LocalMux t4171 (
    .I(seg_12_6_sp4_v_b_5_45515),
    .O(seg_12_6_local_g0_5_49610)
  );
  LocalMux t4172 (
    .I(seg_12_4_lutff_0_out_45487),
    .O(seg_12_4_local_g1_0_49367)
  );
  LocalMux t4173 (
    .I(seg_12_3_neigh_op_top_3_45490),
    .O(seg_12_3_local_g0_3_49239)
  );
  LocalMux t4174 (
    .I(seg_12_4_lutff_4_out_45491),
    .O(seg_12_4_local_g2_4_49379)
  );
  LocalMux t4175 (
    .I(seg_11_4_neigh_op_rgt_5_45492),
    .O(seg_11_4_local_g3_5_45557)
  );
  LocalMux t4176 (
    .I(seg_13_3_neigh_op_tnl_5_45492),
    .O(seg_13_3_local_g2_5_53088)
  );
  LocalMux t4177 (
    .I(seg_3_7_sp4_v_b_19_11916),
    .O(seg_3_7_local_g0_3_15883)
  );
  Span4Mux_v3 t4178 (
    .I(seg_3_4_sp4_h_r_6_15613),
    .O(seg_3_7_sp4_v_b_19_11916)
  );
  Span4Mux_h4 t4179 (
    .I(seg_7_4_sp4_h_r_6_30306),
    .O(seg_3_4_sp4_h_r_6_15613)
  );
  Span4Mux_h4 t4180 (
    .I(seg_11_4_sp4_h_r_3_45627),
    .O(seg_7_4_sp4_h_r_6_30306)
  );
  LocalMux t4181 (
    .I(seg_8_16_sp4_h_r_22_31777),
    .O(seg_8_16_local_g1_6_35525)
  );
  Span4Mux_h3 t4182 (
    .I(seg_11_16_sp4_v_b_6_42917),
    .O(seg_8_16_sp4_h_r_22_31777)
  );
  Span4Mux_v4 t4183 (
    .I(seg_11_12_sp4_v_b_3_42420),
    .O(seg_11_16_sp4_v_b_6_42917)
  );
  Span4Mux_v4 t4184 (
    .I(seg_11_8_sp4_v_b_7_41932),
    .O(seg_11_12_sp4_v_b_3_42420)
  );
  Span4Mux_v4 t4185 (
    .I(seg_11_4_sp4_h_r_7_45631),
    .O(seg_11_8_sp4_v_b_7_41932)
  );
  LocalMux t4186 (
    .I(seg_20_6_sp4_h_r_45_68862),
    .O(seg_20_6_local_g2_5_79641)
  );
  Span4Mux_h3 t4187 (
    .I(seg_17_6_sp4_h_l_40_53537),
    .O(seg_20_6_sp4_h_r_45_68862)
  );
  Span4Mux_h4 t4188 (
    .I(seg_13_6_sp4_v_b_5_49346),
    .O(seg_17_6_sp4_h_l_40_53537)
  );
  LocalMux t4189 (
    .I(seg_12_7_sp4_v_b_1_45634),
    .O(seg_12_7_local_g1_1_49737)
  );
  LocalMux t4190 (
    .I(seg_20_6_sp4_v_b_36_76399),
    .O(seg_20_6_local_g2_4_79640)
  );
  Span4Mux_v1 t4191 (
    .I(seg_20_5_sp4_h_l_45_64908),
    .O(seg_20_6_sp4_v_b_36_76399)
  );
  Span4Mux_h4 t4192 (
    .I(seg_16_5_sp4_h_l_37_49576),
    .O(seg_20_5_sp4_h_l_45_64908)
  );
  LocalMux t4193 (
    .I(seg_20_6_sp4_v_b_46_76409),
    .O(seg_20_6_local_g2_6_79642)
  );
  Span4Mux_v1 t4194 (
    .I(seg_20_5_sp4_h_l_43_64906),
    .O(seg_20_6_sp4_v_b_46_76409)
  );
  Span4Mux_h4 t4195 (
    .I(seg_16_5_sp4_h_l_47_49578),
    .O(seg_20_5_sp4_h_l_43_64906)
  );
  LocalMux t4196 (
    .I(seg_15_6_sp4_h_r_30_53538),
    .O(seg_15_6_local_g2_6_61118)
  );
  Span4Mux_h2 t4197 (
    .I(seg_13_6_sp4_v_b_0_49343),
    .O(seg_15_6_sp4_h_r_30_53538)
  );
  LocalMux t4198 (
    .I(seg_8_16_sp4_v_b_2_31420),
    .O(seg_8_16_local_g0_2_35513)
  );
  Span4Mux_v4 t4199 (
    .I(seg_8_12_sp4_v_b_6_30932),
    .O(seg_8_16_sp4_v_b_2_31420)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t42 (
    .carryinitin(),
    .carryinitout(t41)
  );
  CascadeMux t420 (
    .I(net_31223),
    .O(net_31223_cascademuxed)
  );
  Span4Mux_v4 t4200 (
    .I(seg_8_8_sp4_h_r_6_34629),
    .O(seg_8_12_sp4_v_b_6_30932)
  );
  Span4Mux_h4 t4201 (
    .I(seg_12_8_sp4_v_b_1_45757),
    .O(seg_8_8_sp4_h_r_6_34629)
  );
  LocalMux t4202 (
    .I(seg_12_6_lutff_0_out_45733),
    .O(seg_12_6_local_g3_0_49629)
  );
  LocalMux t4203 (
    .I(seg_12_6_lutff_1_out_45734),
    .O(seg_12_6_local_g3_1_49630)
  );
  LocalMux t4204 (
    .I(seg_12_6_lutff_2_out_45735),
    .O(seg_12_6_local_g2_2_49623)
  );
  LocalMux t4205 (
    .I(seg_12_6_lutff_3_out_45736),
    .O(seg_12_6_local_g0_3_49608)
  );
  LocalMux t4206 (
    .I(seg_12_6_lutff_7_out_45740),
    .O(seg_12_6_local_g3_7_49636)
  );
  LocalMux t4207 (
    .I(seg_0_12_sp12_h_r_0_2614),
    .O(seg_0_12_local_g1_0_2528)
  );
  Span12Mux_h12 t4208 (
    .I(seg_12_12_sp12_v_b_0_48932),
    .O(seg_0_12_sp12_h_r_0_2614)
  );
  LocalMux t4209 (
    .I(seg_0_25_sp4_r_v_b_17_5092),
    .O(seg_0_25_local_g3_1_5346)
  );
  CascadeMux t421 (
    .I(net_31229),
    .O(net_31229_cascademuxed)
  );
  Span4Mux_v3 t4210 (
    .I(seg_1_22_sp4_v_b_8_4205),
    .O(seg_0_25_sp4_r_v_b_17_5092)
  );
  Span4Mux_v4 t4211 (
    .I(seg_1_18_sp4_h_r_8_9382),
    .O(seg_1_22_sp4_v_b_8_4205)
  );
  Span4Mux_h4 t4212 (
    .I(seg_5_18_sp4_h_r_8_24999),
    .O(seg_1_18_sp4_h_r_8_9382)
  );
  Span4Mux_h4 t4213 (
    .I(seg_9_18_sp4_v_b_3_35496),
    .O(seg_5_18_sp4_h_r_8_24999)
  );
  Span4Mux_v4 t4214 (
    .I(seg_9_14_sp4_v_b_7_35008),
    .O(seg_9_18_sp4_v_b_3_35496)
  );
  Span4Mux_v4 t4215 (
    .I(seg_9_10_sp4_v_b_11_34520),
    .O(seg_9_14_sp4_v_b_7_35008)
  );
  Span4Mux_v4 t4216 (
    .I(seg_9_6_sp4_h_r_5_38213),
    .O(seg_9_10_sp4_v_b_11_34520)
  );
  LocalMux t4217 (
    .I(seg_0_12_sp4_v_b_17_2093),
    .O(seg_0_12_local_g1_1_2529)
  );
  Span4Mux_v3 t4218 (
    .I(seg_0_9_sp4_h_r_10_2030),
    .O(seg_0_12_sp4_v_b_17_2093)
  );
  Span4Mux_h4 t4219 (
    .I(seg_4_9_sp4_h_r_10_20053),
    .O(seg_0_9_sp4_h_r_10_2030)
  );
  CascadeMux t422 (
    .I(net_31235),
    .O(net_31235_cascademuxed)
  );
  Span4Mux_h4 t4220 (
    .I(seg_8_9_sp4_h_r_10_34746),
    .O(seg_4_9_sp4_h_r_10_20053)
  );
  Span4Mux_h4 t4221 (
    .I(seg_12_9_sp4_v_b_5_45884),
    .O(seg_8_9_sp4_h_r_10_34746)
  );
  LocalMux t4222 (
    .I(seg_0_12_sp4_v_b_13_2089),
    .O(seg_0_12_local_g1_5_2533)
  );
  Span4Mux_v3 t4223 (
    .I(seg_0_9_sp4_h_r_0_2028),
    .O(seg_0_12_sp4_v_b_13_2089)
  );
  Span4Mux_h4 t4224 (
    .I(seg_4_9_sp4_h_r_0_20051),
    .O(seg_0_9_sp4_h_r_0_2028)
  );
  Span4Mux_h4 t4225 (
    .I(seg_8_9_sp4_h_r_0_34744),
    .O(seg_4_9_sp4_h_r_0_20051)
  );
  Span4Mux_h4 t4226 (
    .I(seg_12_9_sp4_v_b_7_45886),
    .O(seg_8_9_sp4_h_r_0_34744)
  );
  LocalMux t4227 (
    .I(seg_0_25_sp4_v_b_9_4670),
    .O(seg_0_25_local_g1_1_5330)
  );
  Span4Mux_v4 t4228 (
    .I(seg_0_21_sp4_v_b_6_3779),
    .O(seg_0_25_sp4_v_b_9_4670)
  );
  Span4Mux_v4 t4229 (
    .I(seg_0_17_sp4_h_r_0_3712),
    .O(seg_0_21_sp4_v_b_6_3779)
  );
  CascadeMux t423 (
    .I(net_31241),
    .O(net_31241_cascademuxed)
  );
  Span4Mux_h4 t4230 (
    .I(seg_4_17_sp4_h_r_9_21046),
    .O(seg_0_17_sp4_h_r_0_3712)
  );
  Span4Mux_h4 t4231 (
    .I(seg_8_17_sp4_h_r_6_35736),
    .O(seg_4_17_sp4_h_r_9_21046)
  );
  Span4Mux_h4 t4232 (
    .I(seg_12_17_sp4_v_b_6_46871),
    .O(seg_8_17_sp4_h_r_6_35736)
  );
  Span4Mux_v4 t4233 (
    .I(seg_12_13_sp4_v_b_10_46383),
    .O(seg_12_17_sp4_v_b_6_46871)
  );
  Span4Mux_v4 t4234 (
    .I(seg_12_9_sp4_v_b_7_45886),
    .O(seg_12_13_sp4_v_b_10_46383)
  );
  LocalMux t4235 (
    .I(seg_0_25_sp4_v_b_2_4665),
    .O(seg_0_25_local_g1_2_5331)
  );
  Span4Mux_v4 t4236 (
    .I(seg_0_21_sp4_h_r_2_4614),
    .O(seg_0_25_sp4_v_b_2_4665)
  );
  Span4Mux_h4 t4237 (
    .I(seg_4_21_sp4_v_b_9_17347),
    .O(seg_0_21_sp4_h_r_2_4614)
  );
  Span4Mux_v4 t4238 (
    .I(seg_4_17_sp4_h_r_3_21040),
    .O(seg_4_21_sp4_v_b_9_17347)
  );
  Span4Mux_h4 t4239 (
    .I(seg_8_17_sp4_h_r_0_35728),
    .O(seg_4_17_sp4_h_r_3_21040)
  );
  CascadeMux t424 (
    .I(net_31247),
    .O(net_31247_cascademuxed)
  );
  Span4Mux_h4 t4240 (
    .I(seg_12_17_sp4_v_b_0_46865),
    .O(seg_8_17_sp4_h_r_0_35728)
  );
  Span4Mux_v4 t4241 (
    .I(seg_12_13_sp4_v_b_9_46380),
    .O(seg_12_17_sp4_v_b_0_46865)
  );
  Span4Mux_v4 t4242 (
    .I(seg_12_9_sp4_v_b_9_45888),
    .O(seg_12_13_sp4_v_b_9_46380)
  );
  LocalMux t4243 (
    .I(seg_13_7_neigh_op_lft_0_45856),
    .O(seg_13_7_local_g0_0_53559)
  );
  LocalMux t4244 (
    .I(seg_13_6_neigh_op_tnl_1_45857),
    .O(seg_13_6_local_g2_1_53453)
  );
  LocalMux t4245 (
    .I(seg_12_7_lutff_6_out_45862),
    .O(seg_12_7_local_g1_6_49742)
  );
  LocalMux t4246 (
    .I(seg_13_7_neigh_op_lft_7_45863),
    .O(seg_13_7_local_g0_7_53566)
  );
  LocalMux t4247 (
    .I(seg_10_19_sp4_r_v_b_7_43285),
    .O(seg_10_19_local_g1_7_43557)
  );
  Span4Mux_v4 t4248 (
    .I(seg_11_15_sp4_v_b_11_42797),
    .O(seg_10_19_sp4_r_v_b_7_43285)
  );
  Span4Mux_v4 t4249 (
    .I(seg_11_11_sp4_v_b_11_42305),
    .O(seg_11_15_sp4_v_b_11_42797)
  );
  CascadeMux t425 (
    .I(net_31253),
    .O(net_31253_cascademuxed)
  );
  Span4Mux_v4 t4250 (
    .I(seg_11_7_sp4_h_r_11_45994),
    .O(seg_11_11_sp4_v_b_11_42305)
  );
  LocalMux t4251 (
    .I(seg_14_6_sp4_v_b_13_53297),
    .O(seg_14_6_local_g1_5_57279)
  );
  Span4Mux_v1 t4252 (
    .I(seg_14_7_sp4_h_l_37_42160),
    .O(seg_14_6_sp4_v_b_13_53297)
  );
  LocalMux t4253 (
    .I(seg_20_6_sp4_v_b_33_76305),
    .O(seg_20_6_local_g3_1_79645)
  );
  Span4Mux_v2 t4254 (
    .I(seg_20_8_sp4_h_l_38_65272),
    .O(seg_20_6_sp4_v_b_33_76305)
  );
  Span4Mux_h4 t4255 (
    .I(seg_16_8_sp4_h_l_37_49945),
    .O(seg_20_8_sp4_h_l_38_65272)
  );
  LocalMux t4256 (
    .I(seg_20_7_sp4_v_b_22_76307),
    .O(seg_20_7_local_g1_6_79757)
  );
  Span4Mux_v1 t4257 (
    .I(seg_20_8_sp4_h_l_46_65270),
    .O(seg_20_7_sp4_v_b_22_76307)
  );
  Span4Mux_h4 t4258 (
    .I(seg_16_8_sp4_h_l_45_49955),
    .O(seg_20_8_sp4_h_l_46_65270)
  );
  LocalMux t4259 (
    .I(seg_15_6_sp4_h_r_27_53535),
    .O(seg_15_6_local_g2_3_61115)
  );
  CascadeMux t426 (
    .I(net_31259),
    .O(net_31259_cascademuxed)
  );
  Span4Mux_h2 t4260 (
    .I(seg_13_6_sp4_v_t_38_49836),
    .O(seg_15_6_sp4_h_r_27_53535)
  );
  LocalMux t4261 (
    .I(seg_15_18_sp4_r_v_b_12_62432),
    .O(seg_15_18_local_g2_4_62592)
  );
  Span4Mux_v3 t4262 (
    .I(seg_16_15_sp4_v_b_5_61944),
    .O(seg_15_18_sp4_r_v_b_12_62432)
  );
  Span4Mux_v4 t4263 (
    .I(seg_16_11_sp4_h_l_40_50321),
    .O(seg_16_15_sp4_v_b_5_61944)
  );
  Span4Mux_h4 t4264 (
    .I(seg_12_11_sp4_v_b_11_46136),
    .O(seg_16_11_sp4_h_l_40_50321)
  );
  LocalMux t4265 (
    .I(seg_17_8_sp4_r_v_b_18_68870),
    .O(seg_17_8_local_g3_2_69030)
  );
  Span4Mux_v1 t4266 (
    .I(seg_18_9_sp4_h_l_42_57738),
    .O(seg_17_8_sp4_r_v_b_18_68870)
  );
  Span4Mux_h4 t4267 (
    .I(seg_14_9_sp4_h_l_41_42412),
    .O(seg_18_9_sp4_h_l_42_57738)
  );
  LocalMux t4268 (
    .I(seg_17_8_sp4_r_v_b_16_68868),
    .O(seg_17_8_local_g3_0_69028)
  );
  Span4Mux_v1 t4269 (
    .I(seg_18_9_sp4_h_l_46_57732),
    .O(seg_17_8_sp4_r_v_b_16_68868)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t427 (
    .carryinitin(net_35093),
    .carryinitout(net_35137)
  );
  Span4Mux_h4 t4270 (
    .I(seg_14_9_sp4_h_l_45_42416),
    .O(seg_18_9_sp4_h_l_46_57732)
  );
  LocalMux t4271 (
    .I(seg_17_8_sp4_h_r_2_69102),
    .O(seg_17_8_local_g1_2_69014)
  );
  Span4Mux_h0 t4272 (
    .I(seg_17_8_sp4_h_l_43_53784),
    .O(seg_17_8_sp4_h_r_2_69102)
  );
  Span4Mux_h4 t4273 (
    .I(seg_13_8_sp4_v_t_43_50087),
    .O(seg_17_8_sp4_h_l_43_53784)
  );
  LocalMux t4274 (
    .I(seg_11_10_neigh_op_rgt_1_46226),
    .O(seg_11_10_local_g2_1_46283)
  );
  LocalMux t4275 (
    .I(seg_11_14_sp4_v_b_3_42666),
    .O(seg_11_14_local_g0_3_46761)
  );
  Span4Mux_v4 t4276 (
    .I(seg_11_10_sp4_h_r_3_46365),
    .O(seg_11_14_sp4_v_b_3_42666)
  );
  LocalMux t4277 (
    .I(seg_8_10_sp4_h_r_23_31038),
    .O(seg_8_10_local_g1_7_34788)
  );
  Span4Mux_h3 t4278 (
    .I(seg_11_10_sp4_h_r_7_46369),
    .O(seg_8_10_sp4_h_r_23_31038)
  );
  LocalMux t4279 (
    .I(seg_9_14_sp4_v_b_11_35012),
    .O(seg_9_14_local_g1_3_39107)
  );
  CascadeMux t428 (
    .I(net_31364),
    .O(net_31364_cascademuxed)
  );
  Span4Mux_v4 t4280 (
    .I(seg_9_10_sp4_h_r_11_38701),
    .O(seg_9_14_sp4_v_b_11_35012)
  );
  LocalMux t4281 (
    .I(seg_9_12_sp4_h_r_0_38944),
    .O(seg_9_12_local_g1_0_38858)
  );
  Span4Mux_h4 t4282 (
    .I(seg_13_12_sp4_v_b_7_50086),
    .O(seg_9_12_sp4_h_r_0_38944)
  );
  LocalMux t4283 (
    .I(seg_25_11_sp4_v_b_31_95680),
    .O(seg_25_11_local_g2_7_100173)
  );
  Span4Mux_v2 t4284 (
    .I(seg_25_13_sp4_h_l_36_84407),
    .O(seg_25_11_sp4_v_b_31_95680)
  );
  Span4Mux_h4 t4285 (
    .I(seg_21_13_sp4_h_l_40_69720),
    .O(seg_25_13_sp4_h_l_36_84407)
  );
  Span4Mux_h4 t4286 (
    .I(seg_17_13_sp4_h_l_39_54395),
    .O(seg_21_13_sp4_h_l_40_69720)
  );
  Span4Mux_h4 t4287 (
    .I(seg_13_13_sp4_v_b_2_50206),
    .O(seg_17_13_sp4_h_l_39_54395)
  );
  LocalMux t4288 (
    .I(seg_25_12_sp4_v_b_18_95680),
    .O(seg_25_12_local_g1_2_100310)
  );
  Span4Mux_v1 t4289 (
    .I(seg_25_13_sp4_h_l_36_84407),
    .O(seg_25_12_sp4_v_b_18_95680)
  );
  CascadeMux t429 (
    .I(net_31376),
    .O(net_31376_cascademuxed)
  );
  LocalMux t4290 (
    .I(seg_25_11_sp4_v_b_28_95679),
    .O(seg_25_11_local_g2_4_100170)
  );
  Span4Mux_v2 t4291 (
    .I(seg_25_13_sp4_h_l_41_84412),
    .O(seg_25_11_sp4_v_b_28_95679)
  );
  Span4Mux_h4 t4292 (
    .I(seg_21_13_sp4_h_l_41_69719),
    .O(seg_25_13_sp4_h_l_41_84412)
  );
  Span4Mux_h4 t4293 (
    .I(seg_17_13_sp4_h_l_45_54401),
    .O(seg_21_13_sp4_h_l_41_69719)
  );
  Span4Mux_h4 t4294 (
    .I(seg_13_13_sp4_v_b_8_50212),
    .O(seg_17_13_sp4_h_l_45_54401)
  );
  LocalMux t4295 (
    .I(seg_25_12_sp4_v_b_17_95679),
    .O(seg_25_12_local_g1_1_100309)
  );
  Span4Mux_v1 t4296 (
    .I(seg_25_13_sp4_h_l_41_84412),
    .O(seg_25_12_sp4_v_b_17_95679)
  );
  LocalMux t4297 (
    .I(seg_10_13_sp4_h_r_14_39072),
    .O(seg_10_13_local_g0_6_42810)
  );
  Span4Mux_h3 t4298 (
    .I(seg_13_13_sp4_v_b_10_50214),
    .O(seg_10_13_sp4_h_r_14_39072)
  );
  LocalMux t4299 (
    .I(seg_9_15_sp4_h_r_21_35492),
    .O(seg_9_15_local_g0_5_39224)
  );
  CascadeMux t43 (
    .I(net_8707),
    .O(net_8707_cascademuxed)
  );
  CascadeMux t430 (
    .I(net_31382),
    .O(net_31382_cascademuxed)
  );
  Span4Mux_h3 t4300 (
    .I(seg_12_15_sp4_v_b_3_46620),
    .O(seg_9_15_sp4_h_r_21_35492)
  );
  Span4Mux_v4 t4301 (
    .I(seg_12_11_sp4_v_b_7_46132),
    .O(seg_12_15_sp4_v_b_3_46620)
  );
  LocalMux t4302 (
    .I(seg_10_11_sp4_h_r_31_34999),
    .O(seg_10_11_local_g2_7_42581)
  );
  Span4Mux_h2 t4303 (
    .I(seg_12_11_sp4_v_b_7_46132),
    .O(seg_10_11_sp4_h_r_31_34999)
  );
  LocalMux t4304 (
    .I(seg_11_15_sp4_r_v_b_21_46750),
    .O(seg_11_15_local_g3_5_46910)
  );
  Span4Mux_v3 t4305 (
    .I(seg_12_12_sp4_v_b_0_46250),
    .O(seg_11_15_sp4_r_v_b_21_46750)
  );
  LocalMux t4306 (
    .I(seg_12_19_sp4_v_b_22_47243),
    .O(seg_12_19_local_g1_6_51218)
  );
  Span4Mux_v3 t4307 (
    .I(seg_12_16_sp4_v_b_8_46750),
    .O(seg_12_19_sp4_v_b_22_47243)
  );
  Span4Mux_v4 t4308 (
    .I(seg_12_12_sp4_v_b_0_46250),
    .O(seg_12_16_sp4_v_b_8_46750)
  );
  LocalMux t4309 (
    .I(seg_11_17_sp4_r_v_b_1_46864),
    .O(seg_11_17_local_g1_1_47136)
  );
  CascadeMux t431 (
    .I(net_31505),
    .O(net_31505_cascademuxed)
  );
  Span4Mux_v4 t4310 (
    .I(seg_12_13_sp4_v_b_5_46376),
    .O(seg_11_17_sp4_r_v_b_1_46864)
  );
  LocalMux t4311 (
    .I(seg_12_18_sp4_v_b_4_46992),
    .O(seg_12_18_local_g1_4_51093)
  );
  Span4Mux_v4 t4312 (
    .I(seg_12_14_sp4_v_b_4_46500),
    .O(seg_12_18_sp4_v_b_4_46992)
  );
  Span4Mux_v4 t4313 (
    .I(seg_12_10_sp4_v_b_8_46012),
    .O(seg_12_14_sp4_v_b_4_46500)
  );
  LocalMux t4314 (
    .I(seg_16_12_sp4_v_b_41_61945),
    .O(seg_16_12_local_g2_1_65682)
  );
  Span4Mux_v1 t4315 (
    .I(seg_16_11_sp4_h_l_41_50320),
    .O(seg_16_12_sp4_v_b_41_61945)
  );
  LocalMux t4316 (
    .I(seg_13_19_sp4_v_b_20_51072),
    .O(seg_13_19_local_g0_4_55039)
  );
  Span4Mux_v3 t4317 (
    .I(seg_13_16_sp4_v_b_1_50572),
    .O(seg_13_19_sp4_v_b_20_51072)
  );
  Span4Mux_v4 t4318 (
    .I(seg_13_12_sp4_v_b_10_50091),
    .O(seg_13_16_sp4_v_b_1_50572)
  );
  LocalMux t4319 (
    .I(seg_13_18_sp4_v_b_7_50824),
    .O(seg_13_18_local_g0_7_54919)
  );
  CascadeMux t432 (
    .I(net_31511),
    .O(net_31511_cascademuxed)
  );
  Span4Mux_v4 t4320 (
    .I(seg_13_14_sp4_v_b_4_50331),
    .O(seg_13_18_sp4_v_b_7_50824)
  );
  LocalMux t4321 (
    .I(seg_13_18_sp4_v_b_9_50826),
    .O(seg_13_18_local_g0_1_54913)
  );
  Span4Mux_v4 t4322 (
    .I(seg_13_14_sp4_v_b_6_50333),
    .O(seg_13_18_sp4_v_b_9_50826)
  );
  LocalMux t4323 (
    .I(seg_13_18_sp4_v_b_4_50823),
    .O(seg_13_18_local_g0_4_54916)
  );
  Span4Mux_v4 t4324 (
    .I(seg_13_14_sp4_v_b_8_50335),
    .O(seg_13_18_sp4_v_b_4_50823)
  );
  LocalMux t4325 (
    .I(seg_11_12_neigh_op_rgt_0_46471),
    .O(seg_11_12_local_g3_0_46536)
  );
  LocalMux t4326 (
    .I(seg_12_12_lutff_1_out_46472),
    .O(seg_12_12_local_g3_1_50368)
  );
  LocalMux t4327 (
    .I(seg_16_12_sp4_h_r_6_65767),
    .O(seg_16_12_local_g1_6_65679)
  );
  Span4Mux_h0 t4328 (
    .I(seg_16_12_sp4_h_l_43_50445),
    .O(seg_16_12_sp4_h_r_6_65767)
  );
  LocalMux t4329 (
    .I(seg_12_13_lutff_0_out_46594),
    .O(seg_12_13_local_g0_0_50466)
  );
  CascadeMux t433 (
    .I(net_31592),
    .O(net_31592_cascademuxed)
  );
  LocalMux t4330 (
    .I(seg_11_12_neigh_op_tnr_2_46596),
    .O(seg_11_12_local_g2_2_46530)
  );
  LocalMux t4331 (
    .I(seg_12_12_neigh_op_top_2_46596),
    .O(seg_12_12_local_g1_2_50353)
  );
  LocalMux t4332 (
    .I(seg_13_13_neigh_op_lft_2_46596),
    .O(seg_13_13_local_g0_2_54299)
  );
  LocalMux t4333 (
    .I(seg_13_14_neigh_op_bnl_2_46596),
    .O(seg_13_14_local_g3_2_54446)
  );
  LocalMux t4334 (
    .I(seg_12_13_lutff_3_out_46597),
    .O(seg_12_13_local_g1_3_50477)
  );
  LocalMux t4335 (
    .I(seg_12_13_lutff_4_out_46598),
    .O(seg_12_13_local_g3_4_50494)
  );
  LocalMux t4336 (
    .I(seg_12_13_lutff_6_out_46600),
    .O(seg_12_13_local_g0_6_50472)
  );
  LocalMux t4337 (
    .I(seg_10_11_sp4_r_v_b_33_42549),
    .O(seg_10_11_local_g2_1_42575)
  );
  Span4Mux_v2 t4338 (
    .I(seg_11_13_sp4_h_r_9_46740),
    .O(seg_10_11_sp4_r_v_b_33_42549)
  );
  LocalMux t4339 (
    .I(seg_10_15_sp4_r_v_b_27_43035),
    .O(seg_10_15_local_g0_3_43053)
  );
  CascadeMux t434 (
    .I(net_31598),
    .O(net_31598_cascademuxed)
  );
  Span4Mux_v2 t4340 (
    .I(seg_11_13_sp4_h_r_9_46740),
    .O(seg_10_15_sp4_r_v_b_27_43035)
  );
  LocalMux t4341 (
    .I(seg_10_17_sp4_r_v_b_3_43035),
    .O(seg_10_17_local_g1_3_43307)
  );
  Span4Mux_v4 t4342 (
    .I(seg_11_13_sp4_h_r_9_46740),
    .O(seg_10_17_sp4_r_v_b_3_43035)
  );
  LocalMux t4343 (
    .I(seg_11_17_sp4_v_b_3_43035),
    .O(seg_11_17_local_g1_3_47138)
  );
  Span4Mux_v4 t4344 (
    .I(seg_11_13_sp4_h_r_9_46740),
    .O(seg_11_17_sp4_v_b_3_43035)
  );
  LocalMux t4345 (
    .I(seg_9_13_sp4_h_r_1_39068),
    .O(seg_9_13_local_g1_1_38982)
  );
  LocalMux t4346 (
    .I(seg_9_15_sp4_v_b_25_35371),
    .O(seg_9_15_local_g3_1_39244)
  );
  Span4Mux_v2 t4347 (
    .I(seg_9_13_sp4_h_r_1_39068),
    .O(seg_9_15_sp4_v_b_25_35371)
  );
  LocalMux t4348 (
    .I(seg_9_17_sp4_v_b_1_35371),
    .O(seg_9_17_local_g0_1_39466)
  );
  Span4Mux_v4 t4349 (
    .I(seg_9_13_sp4_h_r_1_39068),
    .O(seg_9_17_sp4_v_b_1_35371)
  );
  CascadeMux t435 (
    .I(net_31604),
    .O(net_31604_cascademuxed)
  );
  LocalMux t4350 (
    .I(seg_11_13_sp4_h_r_25_39068),
    .O(seg_11_13_local_g3_1_46660)
  );
  LocalMux t4351 (
    .I(seg_13_15_sp4_v_b_13_50573),
    .O(seg_13_15_local_g1_5_54556)
  );
  LocalMux t4352 (
    .I(seg_14_8_sp4_h_r_21_53786),
    .O(seg_14_8_local_g0_5_57517)
  );
  Span4Mux_h1 t4353 (
    .I(seg_13_8_sp4_v_t_38_50082),
    .O(seg_14_8_sp4_h_r_21_53786)
  );
  Span4Mux_v4 t4354 (
    .I(seg_13_12_sp4_v_t_37_50573),
    .O(seg_13_8_sp4_v_t_38_50082)
  );
  LocalMux t4355 (
    .I(seg_12_15_sp4_r_v_b_19_50579),
    .O(seg_12_15_local_g3_3_50739)
  );
  LocalMux t4356 (
    .I(seg_12_16_sp4_r_v_b_6_50579),
    .O(seg_12_16_local_g1_6_50849)
  );
  LocalMux t4357 (
    .I(seg_13_16_sp4_v_b_6_50579),
    .O(seg_13_16_local_g0_6_54672)
  );
  LocalMux t4358 (
    .I(seg_13_8_sp4_v_b_21_49720),
    .O(seg_13_8_local_g0_5_53687)
  );
  Span4Mux_v1 t4359 (
    .I(seg_13_9_sp4_v_t_40_50207),
    .O(seg_13_8_sp4_v_b_21_49720)
  );
  CascadeMux t436 (
    .I(net_31610),
    .O(net_31610_cascademuxed)
  );
  LocalMux t4360 (
    .I(seg_13_10_sp4_v_b_40_50207),
    .O(seg_13_10_local_g2_0_53944)
  );
  LocalMux t4361 (
    .I(seg_13_10_sp4_v_b_40_50207),
    .O(seg_13_10_local_g3_0_53952)
  );
  LocalMux t4362 (
    .I(seg_13_11_sp4_v_b_29_50207),
    .O(seg_13_11_local_g2_5_54072)
  );
  LocalMux t4363 (
    .I(seg_13_17_sp4_v_b_8_50704),
    .O(seg_13_17_local_g0_0_54789)
  );
  Span4Mux_v4 t4364 (
    .I(seg_13_13_sp4_v_b_5_50207),
    .O(seg_13_17_sp4_v_b_8_50704)
  );
  LocalMux t4365 (
    .I(seg_14_9_sp4_h_r_16_53906),
    .O(seg_14_9_local_g0_0_57635)
  );
  Span4Mux_h1 t4366 (
    .I(seg_13_9_sp4_v_t_40_50207),
    .O(seg_14_9_sp4_h_r_16_53906)
  );
  LocalMux t4367 (
    .I(seg_9_14_sp4_h_r_20_35370),
    .O(seg_9_14_local_g0_4_39100)
  );
  Span4Mux_h3 t4368 (
    .I(seg_12_14_sp4_v_b_9_46503),
    .O(seg_9_14_sp4_h_r_20_35370)
  );
  LocalMux t4369 (
    .I(seg_11_11_sp4_r_v_b_44_46503),
    .O(seg_11_11_local_g3_4_46417)
  );
  CascadeMux t437 (
    .I(net_31616),
    .O(net_31616_cascademuxed)
  );
  LocalMux t4370 (
    .I(seg_11_15_sp4_r_v_b_12_46741),
    .O(seg_11_15_local_g2_4_46901)
  );
  LocalMux t4371 (
    .I(seg_12_16_sp4_v_b_1_46741),
    .O(seg_12_16_local_g1_1_50844)
  );
  LocalMux t4372 (
    .I(seg_12_14_lutff_1_out_46718),
    .O(seg_12_14_local_g3_1_50614)
  );
  LocalMux t4373 (
    .I(seg_12_14_lutff_3_out_46720),
    .O(seg_12_14_local_g3_3_50616)
  );
  LocalMux t4374 (
    .I(seg_12_14_lutff_4_out_46721),
    .O(seg_12_14_local_g3_4_50617)
  );
  LocalMux t4375 (
    .I(seg_12_14_lutff_5_out_46722),
    .O(seg_12_14_local_g1_5_50602)
  );
  LocalMux t4376 (
    .I(seg_13_8_sp4_v_b_37_49958),
    .O(seg_13_8_local_g2_5_53703)
  );
  Span4Mux_v3 t4377 (
    .I(seg_13_11_sp4_v_t_37_50450),
    .O(seg_13_8_sp4_v_b_37_49958)
  );
  LocalMux t4378 (
    .I(seg_11_12_sp4_r_v_b_24_46496),
    .O(seg_11_12_local_g0_0_46512)
  );
  LocalMux t4379 (
    .I(seg_13_14_neigh_op_tnl_0_46840),
    .O(seg_13_14_local_g3_0_54444)
  );
  CascadeMux t438 (
    .I(net_31622),
    .O(net_31622_cascademuxed)
  );
  LocalMux t4380 (
    .I(seg_11_15_neigh_op_rgt_2_46842),
    .O(seg_11_15_local_g2_2_46899)
  );
  LocalMux t4381 (
    .I(seg_11_14_neigh_op_tnr_3_46843),
    .O(seg_11_14_local_g3_3_46785)
  );
  LocalMux t4382 (
    .I(seg_13_15_neigh_op_lft_3_46843),
    .O(seg_13_15_local_g1_3_54554)
  );
  LocalMux t4383 (
    .I(seg_13_15_neigh_op_lft_4_46844),
    .O(seg_13_15_local_g1_4_54555)
  );
  LocalMux t4384 (
    .I(seg_12_16_neigh_op_bot_5_46845),
    .O(seg_12_16_local_g0_5_50840)
  );
  LocalMux t4385 (
    .I(seg_15_14_sp4_r_v_b_19_61947),
    .O(seg_15_14_local_g3_3_62107)
  );
  Span4Mux_v1 t4386 (
    .I(seg_16_15_sp4_h_l_37_50806),
    .O(seg_15_14_sp4_r_v_b_19_61947)
  );
  LocalMux t4387 (
    .I(seg_10_13_sp4_r_v_b_26_42790),
    .O(seg_10_13_local_g0_2_42806)
  );
  Span4Mux_v2 t4388 (
    .I(seg_11_15_sp4_h_r_9_46986),
    .O(seg_10_13_sp4_r_v_b_26_42790)
  );
  LocalMux t4389 (
    .I(seg_11_13_sp4_v_b_26_42790),
    .O(seg_11_13_local_g2_2_46653)
  );
  CascadeMux t439 (
    .I(net_31628),
    .O(net_31628_cascademuxed)
  );
  Span4Mux_v2 t4390 (
    .I(seg_11_15_sp4_h_r_9_46986),
    .O(seg_11_13_sp4_v_b_26_42790)
  );
  LocalMux t4391 (
    .I(seg_14_9_sp4_r_v_b_27_57620),
    .O(seg_14_9_local_g1_3_57646)
  );
  Span4Mux_v2 t4392 (
    .I(seg_15_11_sp4_v_t_38_58112),
    .O(seg_14_9_sp4_r_v_b_27_57620)
  );
  Span4Mux_v4 t4393 (
    .I(seg_15_15_sp4_h_l_44_46986),
    .O(seg_15_11_sp4_v_t_38_58112)
  );
  LocalMux t4394 (
    .I(seg_15_9_sp4_v_b_35_57628),
    .O(seg_15_9_local_g3_3_61492)
  );
  Span4Mux_v2 t4395 (
    .I(seg_15_11_sp4_v_t_46_58120),
    .O(seg_15_9_sp4_v_b_35_57628)
  );
  Span4Mux_v4 t4396 (
    .I(seg_15_15_sp4_h_l_46_46978),
    .O(seg_15_11_sp4_v_t_46_58120)
  );
  LocalMux t4397 (
    .I(seg_13_14_sp4_r_v_b_19_54287),
    .O(seg_13_14_local_g3_3_54447)
  );
  Span4Mux_v1 t4398 (
    .I(seg_14_15_sp4_h_l_43_43152),
    .O(seg_13_14_sp4_r_v_b_19_54287)
  );
  LocalMux t4399 (
    .I(seg_14_11_sp4_v_b_2_53791),
    .O(seg_14_11_local_g0_2_57883)
  );
  CascadeMux t44 (
    .I(net_8719),
    .O(net_8719_cascademuxed)
  );
  CascadeMux t440 (
    .I(net_31634),
    .O(net_31634_cascademuxed)
  );
  Span4Mux_v0 t4400 (
    .I(seg_14_11_sp4_v_t_43_54287),
    .O(seg_14_11_sp4_v_b_2_53791)
  );
  Span4Mux_v4 t4401 (
    .I(seg_14_15_sp4_h_l_43_43152),
    .O(seg_14_11_sp4_v_t_43_54287)
  );
  LocalMux t4402 (
    .I(seg_9_13_sp4_r_v_b_34_38967),
    .O(seg_9_13_local_g2_2_38991)
  );
  Span4Mux_v2 t4403 (
    .I(seg_10_15_sp4_h_r_10_43146),
    .O(seg_9_13_sp4_r_v_b_34_38967)
  );
  LocalMux t4404 (
    .I(seg_9_14_sp4_r_v_b_19_38963),
    .O(seg_9_14_local_g3_3_39123)
  );
  Span4Mux_v1 t4405 (
    .I(seg_10_15_sp4_h_l_43_28143),
    .O(seg_9_14_sp4_r_v_b_19_38963)
  );
  Span4Mux_h0 t4406 (
    .I(seg_10_15_sp4_h_r_10_43146),
    .O(seg_10_15_sp4_h_l_43_28143)
  );
  LocalMux t4407 (
    .I(seg_9_17_sp4_r_v_b_34_39459),
    .O(seg_9_17_local_g2_2_39483)
  );
  Span4Mux_v2 t4408 (
    .I(seg_10_15_sp4_h_r_10_43146),
    .O(seg_9_17_sp4_r_v_b_34_39459)
  );
  LocalMux t4409 (
    .I(seg_10_15_sp4_h_r_18_39322),
    .O(seg_10_15_local_g0_2_43052)
  );
  CascadeMux t441 (
    .I(net_31727),
    .O(net_31727_cascademuxed)
  );
  Span4Mux_h3 t4410 (
    .I(seg_13_15_sp4_h_r_4_54643),
    .O(seg_10_15_sp4_h_r_18_39322)
  );
  Span4Mux_h0 t4411 (
    .I(seg_13_15_sp4_h_l_36_39314),
    .O(seg_13_15_sp4_h_r_4_54643)
  );
  LocalMux t4412 (
    .I(seg_9_15_sp4_h_r_3_39318),
    .O(seg_9_15_local_g1_3_39230)
  );
  LocalMux t4413 (
    .I(seg_20_14_sp4_v_b_19_77018),
    .O(seg_20_14_local_g1_3_80615)
  );
  Span4Mux_v1 t4414 (
    .I(seg_20_15_sp4_h_l_37_66128),
    .O(seg_20_14_sp4_v_b_19_77018)
  );
  Span4Mux_h4 t4415 (
    .I(seg_16_15_sp4_h_l_41_50812),
    .O(seg_20_15_sp4_h_l_37_66128)
  );
  LocalMux t4416 (
    .I(seg_9_12_sp4_h_r_2_38948),
    .O(seg_9_12_local_g0_2_38852)
  );
  Span4Mux_h4 t4417 (
    .I(seg_13_12_sp4_v_t_39_50575),
    .O(seg_9_12_sp4_h_r_2_38948)
  );
  LocalMux t4418 (
    .I(seg_13_10_sp4_v_b_35_50090),
    .O(seg_13_10_local_g3_3_53955)
  );
  Span4Mux_v2 t4419 (
    .I(seg_13_12_sp4_v_t_45_50581),
    .O(seg_13_10_sp4_v_b_35_50090)
  );
  LocalMux t4420 (
    .I(seg_9_16_sp4_h_r_10_39438),
    .O(seg_9_16_local_g0_2_39344)
  );
  Span4Mux_h4 t4421 (
    .I(seg_13_16_sp4_v_b_10_50583),
    .O(seg_9_16_sp4_h_r_10_39438)
  );
  LocalMux t4422 (
    .I(seg_12_19_sp4_r_v_b_19_51071),
    .O(seg_12_19_local_g3_3_51231)
  );
  Span4Mux_v3 t4423 (
    .I(seg_13_16_sp4_v_b_10_50583),
    .O(seg_12_19_sp4_r_v_b_19_51071)
  );
  LocalMux t4424 (
    .I(seg_13_7_sp4_h_r_11_53656),
    .O(seg_13_7_local_g1_3_53570)
  );
  Span4Mux_h0 t4425 (
    .I(seg_13_7_sp4_v_t_43_49964),
    .O(seg_13_7_sp4_h_r_11_53656)
  );
  Span4Mux_v4 t4426 (
    .I(seg_13_11_sp4_v_t_38_50451),
    .O(seg_13_7_sp4_v_t_43_49964)
  );
  LocalMux t4427 (
    .I(seg_10_17_sp4_h_r_18_39568),
    .O(seg_10_17_local_g0_2_43298)
  );
  Span4Mux_h3 t4428 (
    .I(seg_13_17_sp4_v_b_7_50701),
    .O(seg_10_17_sp4_h_r_18_39568)
  );
  LocalMux t4429 (
    .I(seg_13_11_sp4_v_b_27_50205),
    .O(seg_13_11_local_g3_3_54078)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t443 (
    .carryinitin(),
    .carryinitout(t442)
  );
  Span4Mux_v2 t4430 (
    .I(seg_13_13_sp4_v_t_42_50701),
    .O(seg_13_11_sp4_v_b_27_50205)
  );
  LocalMux t4431 (
    .I(seg_13_9_sp4_v_b_35_49967),
    .O(seg_13_9_local_g3_3_53832)
  );
  Span4Mux_v2 t4432 (
    .I(seg_13_11_sp4_h_l_40_38828),
    .O(seg_13_9_sp4_v_b_35_49967)
  );
  Span4Mux_h0 t4433 (
    .I(seg_13_11_sp4_v_t_40_50453),
    .O(seg_13_11_sp4_h_l_40_38828)
  );
  LocalMux t4434 (
    .I(seg_13_13_sp4_v_b_35_50459),
    .O(seg_13_13_local_g3_3_54324)
  );
  Span4Mux_v2 t4435 (
    .I(seg_13_11_sp4_h_r_5_54152),
    .O(seg_13_13_sp4_v_b_35_50459)
  );
  Span4Mux_h0 t4436 (
    .I(seg_13_11_sp4_v_t_40_50453),
    .O(seg_13_11_sp4_h_r_5_54152)
  );
  LocalMux t4437 (
    .I(seg_12_11_sp4_r_v_b_3_49959),
    .O(seg_12_11_local_g1_3_50231)
  );
  Span4Mux_v1 t4438 (
    .I(seg_13_11_sp4_v_t_42_50455),
    .O(seg_12_11_sp4_r_v_b_3_49959)
  );
  LocalMux t4439 (
    .I(seg_8_10_sp4_v_b_26_30928),
    .O(seg_8_10_local_g2_2_34791)
  );
  CascadeMux t444 (
    .I(net_31838),
    .O(net_31838_cascademuxed)
  );
  Span4Mux_v2 t4440 (
    .I(seg_8_12_sp4_h_r_9_35124),
    .O(seg_8_10_sp4_v_b_26_30928)
  );
  Span4Mux_h4 t4441 (
    .I(seg_12_12_sp4_v_t_38_46743),
    .O(seg_8_12_sp4_h_r_9_35124)
  );
  LocalMux t4442 (
    .I(seg_12_9_sp4_v_b_43_46256),
    .O(seg_12_9_local_g3_3_50001)
  );
  Span4Mux_v3 t4443 (
    .I(seg_12_12_sp4_v_t_38_46743),
    .O(seg_12_9_sp4_v_b_43_46256)
  );
  LocalMux t4444 (
    .I(seg_13_12_sp4_h_r_18_50446),
    .O(seg_13_12_local_g0_2_54176)
  );
  Span4Mux_h1 t4445 (
    .I(seg_12_12_sp4_v_t_42_46747),
    .O(seg_13_12_sp4_h_r_18_50446)
  );
  LocalMux t4446 (
    .I(seg_10_11_sp4_h_r_26_34994),
    .O(seg_10_11_local_g2_2_42576)
  );
  Span4Mux_h2 t4447 (
    .I(seg_12_11_sp4_v_t_39_46621),
    .O(seg_10_11_sp4_h_r_26_34994)
  );
  LocalMux t4448 (
    .I(seg_10_16_sp4_h_r_26_35609),
    .O(seg_10_16_local_g2_2_43191)
  );
  Span4Mux_h2 t4449 (
    .I(seg_12_16_sp4_v_b_9_46749),
    .O(seg_10_16_sp4_h_r_26_35609)
  );
  LocalMux t4450 (
    .I(seg_11_10_sp4_r_v_b_33_46257),
    .O(seg_11_10_local_g0_2_46268)
  );
  Span4Mux_v2 t4451 (
    .I(seg_12_12_sp4_v_t_44_46749),
    .O(seg_11_10_sp4_r_v_b_33_46257)
  );
  LocalMux t4452 (
    .I(seg_12_12_sp4_h_r_2_50441),
    .O(seg_12_12_local_g0_2_50345)
  );
  Span4Mux_h0 t4453 (
    .I(seg_12_12_sp4_v_t_44_46749),
    .O(seg_12_12_sp4_h_r_2_50441)
  );
  LocalMux t4454 (
    .I(seg_11_17_sp4_r_v_b_10_46875),
    .O(seg_11_17_local_g2_2_47145)
  );
  LocalMux t4455 (
    .I(seg_10_14_sp4_h_r_35_35362),
    .O(seg_10_14_local_g3_3_42954)
  );
  Span4Mux_h2 t4456 (
    .I(seg_12_14_sp4_v_t_46_46997),
    .O(seg_10_14_sp4_h_r_35_35362)
  );
  LocalMux t4457 (
    .I(seg_12_18_sp4_v_b_11_46997),
    .O(seg_12_18_local_g1_3_51092)
  );
  LocalMux t4458 (
    .I(seg_12_17_neigh_op_bot_0_46963),
    .O(seg_12_17_local_g1_0_50966)
  );
  LocalMux t4459 (
    .I(seg_12_17_neigh_op_bot_1_46964),
    .O(seg_12_17_local_g0_1_50959)
  );
  CascadeMux t446 (
    .I(net_31844),
    .O(net_31844_cascademuxed)
  );
  LocalMux t4460 (
    .I(seg_12_15_neigh_op_top_3_46966),
    .O(seg_12_15_local_g0_3_50715)
  );
  LocalMux t4461 (
    .I(seg_12_15_neigh_op_top_3_46966),
    .O(seg_12_15_local_g1_3_50723)
  );
  LocalMux t4462 (
    .I(seg_12_16_lutff_3_out_46966),
    .O(seg_12_16_local_g1_3_50846)
  );
  LocalMux t4463 (
    .I(seg_12_16_lutff_4_out_46967),
    .O(seg_12_16_local_g1_4_50847)
  );
  LocalMux t4464 (
    .I(seg_13_16_neigh_op_lft_4_46967),
    .O(seg_13_16_local_g0_4_54670)
  );
  LocalMux t4465 (
    .I(seg_12_16_lutff_5_out_46968),
    .O(seg_12_16_local_g1_5_50848)
  );
  LocalMux t4466 (
    .I(seg_12_17_neigh_op_bot_5_46968),
    .O(seg_12_17_local_g1_5_50971)
  );
  LocalMux t4467 (
    .I(seg_12_16_lutff_6_out_46969),
    .O(seg_12_16_local_g2_6_50857)
  );
  LocalMux t4468 (
    .I(seg_12_16_lutff_7_out_46970),
    .O(seg_12_16_local_g0_7_50842)
  );
  LocalMux t4469 (
    .I(seg_5_6_sp12_h_r_11_1346),
    .O(seg_5_6_local_g0_3_23422)
  );
  Span12Mux_h7 t4470 (
    .I(seg_12_6_sp12_v_t_23_49698),
    .O(seg_5_6_sp12_h_r_11_1346)
  );
  LocalMux t4471 (
    .I(seg_12_16_neigh_op_top_1_47087),
    .O(seg_12_16_local_g0_1_50836)
  );
  LocalMux t4472 (
    .I(seg_12_16_neigh_op_top_2_47088),
    .O(seg_12_16_local_g0_2_50837)
  );
  LocalMux t4473 (
    .I(seg_12_16_neigh_op_top_3_47089),
    .O(seg_12_16_local_g0_3_50838)
  );
  LocalMux t4474 (
    .I(seg_12_17_lutff_4_out_47090),
    .O(seg_12_17_local_g2_4_50978)
  );
  LocalMux t4475 (
    .I(seg_12_16_neigh_op_top_6_47092),
    .O(seg_12_16_local_g0_6_50841)
  );
  LocalMux t4476 (
    .I(seg_13_16_neigh_op_tnl_6_47092),
    .O(seg_13_16_local_g3_6_54696)
  );
  LocalMux t4477 (
    .I(seg_13_17_neigh_op_lft_6_47092),
    .O(seg_13_17_local_g1_6_54803)
  );
  LocalMux t4478 (
    .I(seg_12_16_neigh_op_top_7_47093),
    .O(seg_12_16_local_g1_7_50850)
  );
  LocalMux t4479 (
    .I(seg_13_17_neigh_op_lft_7_47093),
    .O(seg_13_17_local_g1_7_54804)
  );
  CascadeMux t448 (
    .I(net_31850),
    .O(net_31850_cascademuxed)
  );
  LocalMux t4480 (
    .I(seg_13_15_sp4_v_b_39_50821),
    .O(seg_13_15_local_g3_7_54574)
  );
  LocalMux t4481 (
    .I(seg_12_15_sp4_v_b_36_46987),
    .O(seg_12_15_local_g3_4_50740)
  );
  LocalMux t4482 (
    .I(seg_12_15_sp4_v_b_38_46989),
    .O(seg_12_15_local_g2_6_50734)
  );
  LocalMux t4483 (
    .I(seg_12_15_sp4_v_b_38_46989),
    .O(seg_12_15_local_g3_6_50742)
  );
  LocalMux t4484 (
    .I(seg_11_18_neigh_op_rgt_2_47211),
    .O(seg_11_18_local_g2_2_47268)
  );
  LocalMux t4485 (
    .I(seg_11_18_neigh_op_rgt_4_47213),
    .O(seg_11_18_local_g3_4_47278)
  );
  LocalMux t4486 (
    .I(seg_11_18_neigh_op_tnr_3_47335),
    .O(seg_11_18_local_g3_3_47277)
  );
  GlobalMux t4487 (
    .I(seg_12_31_local_g1_6_52707_i3),
    .O(seg_1_1_glb_netwk_4_9)
  );
  gio2CtrlBuf t4488 (
    .I(seg_12_31_local_g1_6_52707_i2),
    .O(seg_12_31_local_g1_6_52707_i3)
  );
  ICE_GB t4489 (
    .GLOBALBUFFEROUTPUT(seg_12_31_local_g1_6_52707_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_12_31_local_g1_6_52707_i1)
  );
  IoInMux t4490 (
    .I(seg_12_31_local_g1_6_52707),
    .O(seg_12_31_local_g1_6_52707_i1)
  );
  LocalMux t4491 (
    .I(seg_12_31_span4_horz_r_6_48880),
    .O(seg_12_31_local_g1_6_52707)
  );
  LocalMux t4492 (
    .I(seg_4_2_sp4_r_v_b_3_19049),
    .O(seg_4_2_local_g1_3_19107)
  );
  Span4Mux_v1 t4493 (
    .I(seg_5_2_sp4_h_r_10_23023),
    .O(seg_4_2_sp4_r_v_b_3_19049)
  );
  Span4Mux_h4 t4494 (
    .I(seg_9_2_sp4_h_r_2_37718),
    .O(seg_5_2_sp4_h_r_10_23023)
  );
  Span4Mux_h4 t4495 (
    .I(seg_13_2_sp4_v_b_9_49073),
    .O(seg_9_2_sp4_h_r_2_37718)
  );
  LocalMux t4496 (
    .I(seg_3_1_sp4_h_r_34_6839),
    .O(seg_3_1_local_g2_2_15120)
  );
  Span4Mux_h2 t4497 (
    .I(seg_5_1_sp4_h_r_7_22871),
    .O(seg_3_1_sp4_h_r_34_6839)
  );
  Span4Mux_h4 t4498 (
    .I(seg_9_1_sp4_h_r_4_37561),
    .O(seg_5_1_sp4_h_r_7_22871)
  );
  Span4Mux_h4 t4499 (
    .I(seg_13_1_sp4_v_b_4_49094),
    .O(seg_9_1_sp4_h_r_4_37561)
  );
  CascadeMux t45 (
    .I(net_8743),
    .O(net_8743_cascademuxed)
  );
  CascadeMux t450 (
    .I(net_31856),
    .O(net_31856_cascademuxed)
  );
  LocalMux t4500 (
    .I(seg_13_1_lutff_3_out_48911),
    .O(seg_13_1_local_g1_3_52792)
  );
  LocalMux t4501 (
    .I(seg_13_2_neigh_op_bot_3_48911),
    .O(seg_13_2_local_g1_3_52955)
  );
  LocalMux t4502 (
    .I(seg_14_1_neigh_op_lft_3_48911),
    .O(seg_14_1_local_g0_3_56614)
  );
  GlobalMux t4503 (
    .I(seg_12_0_local_g0_5_48897_i3),
    .O(seg_2_10_glb_netwk_5_10)
  );
  gio2CtrlBuf t4504 (
    .I(seg_12_0_local_g0_5_48897_i2),
    .O(seg_12_0_local_g0_5_48897_i3)
  );
  ICE_GB t4505 (
    .GLOBALBUFFEROUTPUT(seg_12_0_local_g0_5_48897_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_12_0_local_g0_5_48897_i1)
  );
  IoInMux t4506 (
    .I(seg_12_0_local_g0_5_48897),
    .O(seg_12_0_local_g0_5_48897_i1)
  );
  LocalMux t4507 (
    .I(seg_12_0_logic_op_tnr_5_48913),
    .O(seg_12_0_local_g0_5_48897)
  );
  LocalMux t4508 (
    .I(seg_5_17_sp4_v_b_8_20687),
    .O(seg_5_17_local_g0_0_24772)
  );
  Span4Mux_v4 t4509 (
    .I(seg_5_13_sp4_h_r_2_24378),
    .O(seg_5_17_sp4_v_b_8_20687)
  );
  Span4Mux_h4 t4510 (
    .I(seg_9_13_sp4_h_r_6_39075),
    .O(seg_5_13_sp4_h_r_2_24378)
  );
  Span4Mux_h4 t4511 (
    .I(seg_13_13_sp4_v_b_1_50203),
    .O(seg_9_13_sp4_h_r_6_39075)
  );
  Sp12to4 t4512 (
    .I(seg_13_12_sp12_v_b_1_52762),
    .O(seg_13_13_sp4_v_b_1_50203)
  );
  LocalMux t4513 (
    .I(seg_12_13_sp4_r_v_b_1_50203),
    .O(seg_12_13_local_g1_1_50475)
  );
  Sp12to4 t4514 (
    .I(seg_13_12_sp12_v_b_1_52762),
    .O(seg_12_13_sp4_r_v_b_1_50203)
  );
  LocalMux t4515 (
    .I(seg_4_5_sp4_v_b_5_15375),
    .O(seg_4_5_local_g0_5_19470)
  );
  Span4Mux_v4 t4516 (
    .I(seg_4_1_sp4_h_r_5_19038),
    .O(seg_4_5_sp4_v_b_5_15375)
  );
  Span4Mux_h4 t4517 (
    .I(seg_8_1_sp4_h_r_2_33728),
    .O(seg_4_1_sp4_h_r_5_19038)
  );
  Span4Mux_h4 t4518 (
    .I(seg_12_1_sp4_h_r_11_49051),
    .O(seg_8_1_sp4_h_r_2_33728)
  );
  LocalMux t4519 (
    .I(seg_16_3_sp4_v_b_28_60715),
    .O(seg_16_3_local_g3_4_64586)
  );
  CascadeMux t452 (
    .I(net_31862),
    .O(net_31862_cascademuxed)
  );
  Span4Mux_v2 t4520 (
    .I(seg_16_1_sp4_h_l_46_49051),
    .O(seg_16_3_sp4_v_b_28_60715)
  );
  GlobalMux t4521 (
    .I(seg_6_31_local_g0_1_29708_i3),
    .O(seg_2_7_glb_netwk_3_8)
  );
  gio2CtrlBuf t4522 (
    .I(seg_6_31_local_g0_1_29708_i2),
    .O(seg_6_31_local_g0_1_29708_i3)
  );
  ICE_GB t4523 (
    .GLOBALBUFFEROUTPUT(seg_6_31_local_g0_1_29708_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_6_31_local_g0_1_29708_i1)
  );
  IoInMux t4524 (
    .I(seg_6_31_local_g0_1_29708),
    .O(seg_6_31_local_g0_1_29708_i1)
  );
  LocalMux t4525 (
    .I(seg_6_31_span4_vert_33_26481),
    .O(seg_6_31_local_g0_1_29708)
  );
  Span4Mux_v2 t4526 (
    .I(seg_6_29_sp4_h_r_3_29568),
    .O(seg_6_31_span4_vert_33_26481)
  );
  Span4Mux_h4 t4527 (
    .I(seg_10_29_sp4_v_b_3_40680),
    .O(seg_6_29_sp4_h_r_3_29568)
  );
  Span4Mux_v4 t4528 (
    .I(seg_10_25_sp4_v_b_7_40192),
    .O(seg_10_29_sp4_v_b_3_40680)
  );
  Span4Mux_v4 t4529 (
    .I(seg_10_21_sp4_v_b_7_39700),
    .O(seg_10_25_sp4_v_b_7_40192)
  );
  Span4Mux_v4 t4530 (
    .I(seg_10_17_sp4_v_b_4_39207),
    .O(seg_10_21_sp4_v_b_7_39700)
  );
  Span4Mux_v4 t4531 (
    .I(seg_10_13_sp4_v_b_1_38710),
    .O(seg_10_17_sp4_v_b_4_39207)
  );
  Span4Mux_v4 t4532 (
    .I(seg_10_9_sp4_v_b_5_38222),
    .O(seg_10_13_sp4_v_b_1_38710)
  );
  Span4Mux_v4 t4533 (
    .I(seg_10_5_sp4_v_b_9_37734),
    .O(seg_10_9_sp4_v_b_5_38222)
  );
  Span4Mux_v4 t4534 (
    .I(seg_10_1_sp4_h_r_9_41397),
    .O(seg_10_5_sp4_v_b_9_37734)
  );
  LocalMux t4535 (
    .I(seg_4_7_sp4_r_v_b_16_19575),
    .O(seg_4_7_local_g3_0_19735)
  );
  Span4Mux_v3 t4536 (
    .I(seg_5_4_sp4_h_r_11_23270),
    .O(seg_4_7_sp4_r_v_b_16_19575)
  );
  Span4Mux_h4 t4537 (
    .I(seg_9_4_sp4_h_r_3_37965),
    .O(seg_5_4_sp4_h_r_11_23270)
  );
  Span4Mux_h4 t4538 (
    .I(seg_13_4_sp4_v_b_3_49092),
    .O(seg_9_4_sp4_h_r_3_37965)
  );
  LocalMux t4539 (
    .I(seg_13_4_sp4_v_b_3_49092),
    .O(seg_13_4_local_g1_3_53201)
  );
  CascadeMux t454 (
    .I(net_31868),
    .O(net_31868_cascademuxed)
  );
  LocalMux t4540 (
    .I(seg_13_2_lutff_0_out_49036),
    .O(seg_13_2_local_g1_0_52952)
  );
  LocalMux t4541 (
    .I(seg_14_1_neigh_op_tnl_0_49036),
    .O(seg_14_1_local_g2_0_56627)
  );
  LocalMux t4542 (
    .I(seg_12_1_neigh_op_tnr_1_49037),
    .O(seg_12_1_local_g2_1_48967)
  );
  LocalMux t4543 (
    .I(seg_12_1_neigh_op_tnr_1_49037),
    .O(seg_12_1_local_g3_1_48975)
  );
  LocalMux t4544 (
    .I(seg_13_1_neigh_op_top_2_49038),
    .O(seg_13_1_local_g1_2_52791)
  );
  LocalMux t4545 (
    .I(seg_13_2_lutff_2_out_49038),
    .O(seg_13_2_local_g1_2_52954)
  );
  LocalMux t4546 (
    .I(seg_13_1_neigh_op_top_3_49039),
    .O(seg_13_1_local_g0_3_52784)
  );
  LocalMux t4547 (
    .I(seg_13_2_lutff_3_out_49039),
    .O(seg_13_2_local_g2_3_52963)
  );
  LocalMux t4548 (
    .I(seg_13_1_neigh_op_top_4_49040),
    .O(seg_13_1_local_g0_4_52785)
  );
  LocalMux t4549 (
    .I(seg_13_2_lutff_4_out_49040),
    .O(seg_13_2_local_g0_4_52948)
  );
  LocalMux t4550 (
    .I(seg_13_4_sp4_r_v_b_1_52921),
    .O(seg_13_4_local_g1_1_53199)
  );
  LocalMux t4551 (
    .I(seg_13_4_sp4_r_v_b_13_53051),
    .O(seg_13_4_local_g2_5_53211)
  );
  LocalMux t4552 (
    .I(seg_13_3_lutff_0_out_49195),
    .O(seg_13_3_local_g2_0_53083)
  );
  LocalMux t4553 (
    .I(seg_14_4_neigh_op_bnl_1_49196),
    .O(seg_14_4_local_g3_1_57045)
  );
  LocalMux t4554 (
    .I(seg_12_2_neigh_op_tnr_2_49197),
    .O(seg_12_2_local_g2_2_49131)
  );
  LocalMux t4555 (
    .I(seg_13_3_lutff_4_out_49199),
    .O(seg_13_3_local_g2_4_53087)
  );
  LocalMux t4556 (
    .I(seg_12_3_neigh_op_rgt_6_49201),
    .O(seg_12_3_local_g2_6_49258)
  );
  LocalMux t4557 (
    .I(seg_13_2_neigh_op_top_7_49202),
    .O(seg_13_2_local_g1_7_52959)
  );
  LocalMux t4558 (
    .I(seg_25_6_sp4_v_b_19_94847),
    .O(seg_25_6_local_g0_3_99373)
  );
  Span4Mux_v3 t4559 (
    .I(seg_25_3_sp4_h_l_36_83177),
    .O(seg_25_6_sp4_v_b_19_94847)
  );
  CascadeMux t456 (
    .I(net_31874),
    .O(net_31874_cascademuxed)
  );
  Span4Mux_h4 t4560 (
    .I(seg_21_3_sp4_h_l_36_68484),
    .O(seg_25_3_sp4_h_l_36_83177)
  );
  Span4Mux_h4 t4561 (
    .I(seg_17_3_sp4_h_l_47_53163),
    .O(seg_21_3_sp4_h_l_36_68484)
  );
  LocalMux t4562 (
    .I(seg_25_7_sp4_v_b_6_94847),
    .O(seg_25_7_local_g1_6_99534)
  );
  Span4Mux_v4 t4563 (
    .I(seg_25_3_sp4_h_l_36_83177),
    .O(seg_25_7_sp4_v_b_6_94847)
  );
  LocalMux t4564 (
    .I(seg_13_6_sp4_v_b_21_49474),
    .O(seg_13_6_local_g0_5_53441)
  );
  Span4Mux_v3 t4565 (
    .I(seg_13_3_sp4_h_r_2_53165),
    .O(seg_13_6_sp4_v_b_21_49474)
  );
  LocalMux t4566 (
    .I(seg_17_2_sp4_v_b_15_64401),
    .O(seg_17_2_local_g1_7_68281)
  );
  Span4Mux_v1 t4567 (
    .I(seg_17_3_sp4_h_l_39_53165),
    .O(seg_17_2_sp4_v_b_15_64401)
  );
  LocalMux t4568 (
    .I(seg_15_5_sp4_h_r_16_57244),
    .O(seg_15_5_local_g0_0_60973)
  );
  Span4Mux_h1 t4569 (
    .I(seg_14_5_sp4_v_b_11_53060),
    .O(seg_15_5_sp4_h_r_16_57244)
  );
  CascadeMux t457 (
    .I(net_31961),
    .O(net_31961_cascademuxed)
  );
  LocalMux t4570 (
    .I(seg_13_5_sp4_v_b_10_49230),
    .O(seg_13_5_local_g0_2_53315)
  );
  LocalMux t4571 (
    .I(seg_12_4_neigh_op_rgt_0_49318),
    .O(seg_12_4_local_g3_0_49383)
  );
  LocalMux t4572 (
    .I(seg_14_4_neigh_op_lft_0_49318),
    .O(seg_14_4_local_g0_0_57020)
  );
  LocalMux t4573 (
    .I(seg_12_4_neigh_op_rgt_3_49321),
    .O(seg_12_4_local_g3_3_49386)
  );
  LocalMux t4574 (
    .I(seg_13_5_neigh_op_bot_3_49321),
    .O(seg_13_5_local_g1_3_53324)
  );
  LocalMux t4575 (
    .I(seg_14_5_neigh_op_bnl_3_49321),
    .O(seg_14_5_local_g3_3_57170)
  );
  LocalMux t4576 (
    .I(seg_12_5_neigh_op_bnr_4_49322),
    .O(seg_12_5_local_g1_4_49494)
  );
  LocalMux t4577 (
    .I(seg_14_5_neigh_op_bnl_4_49322),
    .O(seg_14_5_local_g2_4_57163)
  );
  LocalMux t4578 (
    .I(seg_13_4_lutff_5_out_49323),
    .O(seg_13_4_local_g1_5_53203)
  );
  LocalMux t4579 (
    .I(seg_12_3_neigh_op_tnr_6_49324),
    .O(seg_12_3_local_g3_6_49266)
  );
  CascadeMux t458 (
    .I(net_31979),
    .O(net_31979_cascademuxed)
  );
  LocalMux t4580 (
    .I(seg_8_6_sp4_v_b_35_30443),
    .O(seg_8_6_local_g2_3_34300)
  );
  Span4Mux_v2 t4581 (
    .I(seg_8_4_sp4_h_r_5_34136),
    .O(seg_8_6_sp4_v_b_35_30443)
  );
  Span4Mux_h4 t4582 (
    .I(seg_12_4_sp4_h_r_5_49460),
    .O(seg_8_4_sp4_h_r_5_34136)
  );
  LocalMux t4583 (
    .I(seg_8_7_sp4_v_b_22_30443),
    .O(seg_8_7_local_g1_6_34418)
  );
  Span4Mux_v3 t4584 (
    .I(seg_8_4_sp4_h_r_5_34136),
    .O(seg_8_7_sp4_v_b_22_30443)
  );
  LocalMux t4585 (
    .I(seg_15_4_sp4_h_r_40_49460),
    .O(seg_15_4_local_g3_0_60874)
  );
  LocalMux t4586 (
    .I(seg_8_6_sp4_v_b_33_30441),
    .O(seg_8_6_local_g3_1_34306)
  );
  Span4Mux_v2 t4587 (
    .I(seg_8_4_sp4_h_r_9_34140),
    .O(seg_8_6_sp4_v_b_33_30441)
  );
  Span4Mux_h4 t4588 (
    .I(seg_12_4_sp4_h_r_9_49464),
    .O(seg_8_4_sp4_h_r_9_34140)
  );
  LocalMux t4589 (
    .I(seg_9_4_sp4_h_r_20_34140),
    .O(seg_9_4_local_g0_4_37870)
  );
  CascadeMux t459 (
    .I(net_31991),
    .O(net_31991_cascademuxed)
  );
  Span4Mux_h3 t4590 (
    .I(seg_12_4_sp4_h_r_9_49464),
    .O(seg_9_4_sp4_h_r_20_34140)
  );
  LocalMux t4591 (
    .I(seg_3_6_sp4_r_v_b_34_15751),
    .O(seg_3_6_local_g2_2_15775)
  );
  Span4Mux_v2 t4592 (
    .I(seg_4_4_sp4_h_r_10_19438),
    .O(seg_3_6_sp4_r_v_b_34_15751)
  );
  Span4Mux_h4 t4593 (
    .I(seg_8_4_sp4_h_r_2_34133),
    .O(seg_4_4_sp4_h_r_10_19438)
  );
  Span4Mux_h4 t4594 (
    .I(seg_12_4_sp4_h_r_11_49456),
    .O(seg_8_4_sp4_h_r_2_34133)
  );
  LocalMux t4595 (
    .I(seg_8_3_sp4_v_b_18_29942),
    .O(seg_8_3_local_g0_2_33914)
  );
  Span4Mux_v1 t4596 (
    .I(seg_8_4_sp4_h_r_2_34133),
    .O(seg_8_3_sp4_v_b_18_29942)
  );
  LocalMux t4597 (
    .I(seg_9_4_sp4_h_r_18_34138),
    .O(seg_9_4_local_g0_2_37868)
  );
  Span4Mux_h3 t4598 (
    .I(seg_12_4_sp4_h_r_11_49456),
    .O(seg_9_4_sp4_h_r_18_34138)
  );
  LocalMux t4599 (
    .I(seg_10_4_sp4_h_r_1_41792),
    .O(seg_10_4_local_g1_1_41706)
  );
  CascadeMux t460 (
    .I(net_32084),
    .O(net_32084_cascademuxed)
  );
  LocalMux t4600 (
    .I(seg_10_6_sp4_v_b_25_38095),
    .O(seg_10_6_local_g2_1_41960)
  );
  Span4Mux_v2 t4601 (
    .I(seg_10_4_sp4_h_r_1_41792),
    .O(seg_10_6_sp4_v_b_25_38095)
  );
  LocalMux t4602 (
    .I(seg_2_8_sp4_h_r_2_12270),
    .O(seg_2_8_local_g0_2_12174)
  );
  Span4Mux_h4 t4603 (
    .I(seg_6_8_sp4_v_b_9_23410),
    .O(seg_2_8_sp4_h_r_2_12270)
  );
  Span4Mux_v4 t4604 (
    .I(seg_6_4_sp4_h_r_3_27018),
    .O(seg_6_8_sp4_v_b_9_23410)
  );
  Span4Mux_h4 t4605 (
    .I(seg_10_4_sp4_h_r_3_41796),
    .O(seg_6_4_sp4_h_r_3_27018)
  );
  LocalMux t4606 (
    .I(seg_5_3_sp4_r_v_b_19_22912),
    .O(seg_5_3_local_g3_3_23077)
  );
  Span4Mux_v1 t4607 (
    .I(seg_6_4_sp4_h_r_6_27021),
    .O(seg_5_3_sp4_r_v_b_19_22912)
  );
  Span4Mux_h4 t4608 (
    .I(seg_10_4_sp4_h_r_3_41796),
    .O(seg_6_4_sp4_h_r_6_27021)
  );
  LocalMux t4609 (
    .I(seg_10_12_sp4_v_b_3_38589),
    .O(seg_10_12_local_g1_3_42692)
  );
  CascadeMux t461 (
    .I(net_32102),
    .O(net_32102_cascademuxed)
  );
  Span4Mux_v4 t4610 (
    .I(seg_10_8_sp4_v_b_3_38097),
    .O(seg_10_12_sp4_v_b_3_38589)
  );
  Span4Mux_v4 t4611 (
    .I(seg_10_4_sp4_h_r_3_41796),
    .O(seg_10_8_sp4_v_b_3_38097)
  );
  LocalMux t4612 (
    .I(seg_15_4_sp4_h_r_28_53290),
    .O(seg_15_4_local_g3_4_60878)
  );
  LocalMux t4613 (
    .I(seg_15_4_sp4_h_r_32_53294),
    .O(seg_15_4_local_g2_0_60866)
  );
  LocalMux t4614 (
    .I(seg_11_5_sp4_h_r_18_41923),
    .O(seg_11_5_local_g0_2_45653)
  );
  Span4Mux_h3 t4615 (
    .I(seg_14_5_sp4_v_b_2_53053),
    .O(seg_11_5_sp4_h_r_18_41923)
  );
  LocalMux t4616 (
    .I(seg_11_2_sp4_h_r_22_41548),
    .O(seg_11_2_local_g1_6_45296)
  );
  Span4Mux_h3 t4617 (
    .I(seg_14_2_sp4_v_t_46_53183),
    .O(seg_11_2_sp4_h_r_22_41548)
  );
  LocalMux t4618 (
    .I(seg_11_7_sp4_h_r_20_42171),
    .O(seg_11_7_local_g1_4_45909)
  );
  Span4Mux_h3 t4619 (
    .I(seg_14_7_sp4_v_b_4_53301),
    .O(seg_11_7_sp4_h_r_20_42171)
  );
  CascadeMux t462 (
    .I(net_33673),
    .O(net_33673_cascademuxed)
  );
  LocalMux t4620 (
    .I(seg_1_7_sp4_h_r_11_7758),
    .O(seg_1_7_local_g1_3_7648)
  );
  Span4Mux_h4 t4621 (
    .I(seg_5_7_sp4_h_r_11_23639),
    .O(seg_1_7_sp4_h_r_11_7758)
  );
  Span4Mux_h4 t4622 (
    .I(seg_9_7_sp4_h_r_3_38334),
    .O(seg_5_7_sp4_h_r_11_23639)
  );
  Span4Mux_h4 t4623 (
    .I(seg_13_7_sp4_v_b_3_49467),
    .O(seg_9_7_sp4_h_r_3_38334)
  );
  LocalMux t4624 (
    .I(seg_9_3_sp4_h_r_3_37842),
    .O(seg_9_3_local_g1_3_37754)
  );
  Span4Mux_h4 t4625 (
    .I(seg_13_3_sp4_v_t_38_49467),
    .O(seg_9_3_sp4_h_r_3_37842)
  );
  LocalMux t4626 (
    .I(seg_12_7_sp4_r_v_b_5_49469),
    .O(seg_12_7_local_g1_5_49741)
  );
  LocalMux t4627 (
    .I(seg_14_6_neigh_op_bnl_0_49441),
    .O(seg_14_6_local_g3_0_57290)
  );
  LocalMux t4628 (
    .I(seg_13_6_neigh_op_bot_1_49442),
    .O(seg_13_6_local_g1_1_53445)
  );
  LocalMux t4629 (
    .I(seg_13_7_sp4_r_v_b_21_53428),
    .O(seg_13_7_local_g3_5_53588)
  );
  CascadeMux t463 (
    .I(net_33824),
    .O(net_33824_cascademuxed)
  );
  LocalMux t4630 (
    .I(seg_13_7_sp4_v_b_2_49468),
    .O(seg_13_7_local_g1_2_53569)
  );
  LocalMux t4631 (
    .I(seg_20_6_sp4_h_r_37_68852),
    .O(seg_20_6_local_g3_5_79649)
  );
  Span4Mux_h3 t4632 (
    .I(seg_17_6_sp4_h_l_37_53530),
    .O(seg_20_6_sp4_h_r_37_68852)
  );
  LocalMux t4633 (
    .I(seg_20_7_sp4_r_v_b_43_79856),
    .O(seg_20_7_local_g3_3_79770)
  );
  Span4Mux_v1 t4634 (
    .I(seg_21_6_sp4_h_l_36_68853),
    .O(seg_20_7_sp4_r_v_b_43_79856)
  );
  Span4Mux_h4 t4635 (
    .I(seg_17_6_sp4_h_l_47_53532),
    .O(seg_21_6_sp4_h_l_36_68853)
  );
  LocalMux t4636 (
    .I(seg_15_6_sp4_h_r_26_53534),
    .O(seg_15_6_local_g2_2_61114)
  );
  LocalMux t4637 (
    .I(seg_15_6_sp4_h_r_44_49710),
    .O(seg_15_6_local_g2_4_61116)
  );
  LocalMux t4638 (
    .I(seg_15_18_sp4_v_b_2_58482),
    .O(seg_15_18_local_g1_2_62582)
  );
  Span4Mux_v4 t4639 (
    .I(seg_15_14_sp4_v_b_11_57997),
    .O(seg_15_18_sp4_v_b_2_58482)
  );
  CascadeMux t464 (
    .I(net_33947),
    .O(net_33947_cascademuxed)
  );
  Span4Mux_v4 t4640 (
    .I(seg_15_10_sp4_v_b_11_57505),
    .O(seg_15_14_sp4_v_b_11_57997)
  );
  Span4Mux_v4 t4641 (
    .I(seg_15_6_sp4_h_l_43_45876),
    .O(seg_15_10_sp4_v_b_11_57505)
  );
  LocalMux t4642 (
    .I(seg_15_6_sp4_h_r_20_57371),
    .O(seg_15_6_local_g1_4_61108)
  );
  Span4Mux_h1 t4643 (
    .I(seg_14_6_sp4_h_l_44_42048),
    .O(seg_15_6_sp4_h_r_20_57371)
  );
  LocalMux t4644 (
    .I(seg_15_6_sp4_h_r_32_53540),
    .O(seg_15_6_local_g2_0_61112)
  );
  LocalMux t4645 (
    .I(seg_15_6_sp4_h_r_12_57361),
    .O(seg_15_6_local_g0_4_61100)
  );
  Span4Mux_h1 t4646 (
    .I(seg_14_6_sp4_v_b_7_53179),
    .O(seg_15_6_sp4_h_r_12_57361)
  );
  LocalMux t4647 (
    .I(seg_14_8_neigh_op_bnl_0_49687),
    .O(seg_14_8_local_g3_0_57536)
  );
  LocalMux t4648 (
    .I(seg_13_8_neigh_op_bot_3_49690),
    .O(seg_13_8_local_g1_3_53693)
  );
  LocalMux t4649 (
    .I(seg_13_8_neigh_op_bot_6_49693),
    .O(seg_13_8_local_g0_6_53688)
  );
  CascadeMux t465 (
    .I(net_33983),
    .O(net_33983_cascademuxed)
  );
  LocalMux t4650 (
    .I(seg_20_7_sp4_h_r_9_79848),
    .O(seg_20_7_local_g1_1_79752)
  );
  Span4Mux_h0 t4651 (
    .I(seg_20_7_sp4_h_l_43_65152),
    .O(seg_20_7_sp4_h_r_9_79848)
  );
  Span4Mux_h4 t4652 (
    .I(seg_16_7_sp4_h_l_38_49827),
    .O(seg_20_7_sp4_h_l_43_65152)
  );
  LocalMux t4653 (
    .I(seg_13_10_sp4_v_b_21_49966),
    .O(seg_13_10_local_g1_5_53941)
  );
  Span4Mux_v3 t4654 (
    .I(seg_13_7_sp4_h_r_2_53657),
    .O(seg_13_10_sp4_v_b_21_49966)
  );
  LocalMux t4655 (
    .I(seg_15_18_sp4_h_r_19_58844),
    .O(seg_15_18_local_g0_3_62575)
  );
  Span4Mux_h1 t4656 (
    .I(seg_14_18_sp4_v_b_0_54650),
    .O(seg_15_18_sp4_h_r_19_58844)
  );
  Span4Mux_v4 t4657 (
    .I(seg_14_14_sp4_v_b_0_54158),
    .O(seg_14_18_sp4_v_b_0_54650)
  );
  Span4Mux_v4 t4658 (
    .I(seg_14_10_sp4_v_b_0_53666),
    .O(seg_14_14_sp4_v_b_0_54158)
  );
  LocalMux t4659 (
    .I(seg_14_9_sp4_v_b_17_53670),
    .O(seg_14_9_local_g0_1_57636)
  );
  CascadeMux t466 (
    .I(net_34205),
    .O(net_34205_cascademuxed)
  );
  LocalMux t4660 (
    .I(seg_13_10_sp4_r_v_b_6_53672),
    .O(seg_13_10_local_g1_6_53942)
  );
  LocalMux t4661 (
    .I(seg_13_8_lutff_5_out_49815),
    .O(seg_13_8_local_g3_5_53711)
  );
  LocalMux t4662 (
    .I(seg_13_8_lutff_6_out_49816),
    .O(seg_13_8_local_g1_6_53696)
  );
  LocalMux t4663 (
    .I(seg_17_8_sp4_h_r_5_69105),
    .O(seg_17_8_local_g0_5_69009)
  );
  Span4Mux_h0 t4664 (
    .I(seg_17_8_sp4_h_l_39_53780),
    .O(seg_17_8_sp4_h_r_5_69105)
  );
  LocalMux t4665 (
    .I(seg_11_12_sp4_r_v_b_3_46251),
    .O(seg_11_12_local_g1_3_46523)
  );
  Span4Mux_v4 t4666 (
    .I(seg_12_8_sp4_h_r_9_49956),
    .O(seg_11_12_sp4_r_v_b_3_46251)
  );
  LocalMux t4667 (
    .I(seg_11_12_sp4_v_b_6_42425),
    .O(seg_11_12_local_g0_6_46518)
  );
  Span4Mux_v4 t4668 (
    .I(seg_11_8_sp4_h_r_0_46114),
    .O(seg_11_12_sp4_v_b_6_42425)
  );
  LocalMux t4669 (
    .I(seg_17_8_sp4_h_r_32_61446),
    .O(seg_17_8_local_g2_0_69020)
  );
  CascadeMux t467 (
    .I(net_34217),
    .O(net_34217_cascademuxed)
  );
  Span4Mux_h2 t4670 (
    .I(seg_15_8_sp4_h_l_45_46124),
    .O(seg_17_8_sp4_h_r_32_61446)
  );
  LocalMux t4671 (
    .I(seg_12_14_sp4_r_v_b_2_50329),
    .O(seg_12_14_local_g1_2_50599)
  );
  Span4Mux_v4 t4672 (
    .I(seg_13_10_sp4_v_b_6_49841),
    .O(seg_12_14_sp4_r_v_b_2_50329)
  );
  LocalMux t4673 (
    .I(seg_13_8_neigh_op_top_2_49935),
    .O(seg_13_8_local_g0_2_53684)
  );
  LocalMux t4674 (
    .I(seg_13_8_neigh_op_top_5_49938),
    .O(seg_13_8_local_g1_5_53695)
  );
  LocalMux t4675 (
    .I(seg_13_10_lutff_1_out_50057),
    .O(seg_13_10_local_g3_1_53953)
  );
  LocalMux t4676 (
    .I(seg_13_10_lutff_2_out_50058),
    .O(seg_13_10_local_g2_2_53946)
  );
  LocalMux t4677 (
    .I(seg_13_11_neigh_op_bot_5_50061),
    .O(seg_13_11_local_g0_5_54056)
  );
  LocalMux t4678 (
    .I(seg_13_18_sp12_v_b_0_53529),
    .O(seg_13_18_local_g3_0_54936)
  );
  LocalMux t4679 (
    .I(seg_16_12_sp4_h_r_25_58099),
    .O(seg_16_12_local_g3_1_65690)
  );
  CascadeMux t468 (
    .I(net_34235),
    .O(net_34235_cascademuxed)
  );
  Span4Mux_h2 t4680 (
    .I(seg_14_12_sp4_v_b_1_53911),
    .O(seg_16_12_sp4_h_r_25_58099)
  );
  LocalMux t4681 (
    .I(seg_13_18_sp12_v_b_5_53774),
    .O(seg_13_18_local_g2_5_54933)
  );
  LocalMux t4682 (
    .I(seg_13_18_sp12_v_b_7_53898),
    .O(seg_13_18_local_g2_7_54935)
  );
  LocalMux t4683 (
    .I(seg_16_12_sp4_r_v_b_45_65780),
    .O(seg_16_12_local_g3_5_65694)
  );
  Span4Mux_v1 t4684 (
    .I(seg_17_11_sp4_h_l_45_54155),
    .O(seg_16_12_sp4_r_v_b_45_65780)
  );
  LocalMux t4685 (
    .I(seg_13_19_sp4_v_b_9_50949),
    .O(seg_13_19_local_g0_1_55036)
  );
  Span4Mux_v4 t4686 (
    .I(seg_13_15_sp4_v_b_1_50449),
    .O(seg_13_19_sp4_v_b_9_50949)
  );
  Span4Mux_v4 t4687 (
    .I(seg_13_11_sp4_v_b_10_49968),
    .O(seg_13_15_sp4_v_b_1_50449)
  );
  LocalMux t4688 (
    .I(seg_13_18_sp4_v_b_5_50822),
    .O(seg_13_18_local_g0_5_54917)
  );
  Span4Mux_v4 t4689 (
    .I(seg_13_14_sp4_v_b_9_50334),
    .O(seg_13_18_sp4_v_b_5_50822)
  );
  CascadeMux t469 (
    .I(net_34346),
    .O(net_34346_cascademuxed)
  );
  LocalMux t4690 (
    .I(seg_13_13_neigh_op_bot_0_50302),
    .O(seg_13_13_local_g1_0_54305)
  );
  LocalMux t4691 (
    .I(seg_13_13_neigh_op_bot_2_50304),
    .O(seg_13_13_local_g1_2_54307)
  );
  LocalMux t4692 (
    .I(seg_13_13_neigh_op_bot_3_50305),
    .O(seg_13_13_local_g1_3_54308)
  );
  LocalMux t4693 (
    .I(seg_13_11_neigh_op_top_4_50306),
    .O(seg_13_11_local_g0_4_54055)
  );
  LocalMux t4694 (
    .I(seg_12_12_neigh_op_rgt_5_50307),
    .O(seg_12_12_local_g3_5_50372)
  );
  LocalMux t4695 (
    .I(seg_13_13_neigh_op_bot_6_50308),
    .O(seg_13_13_local_g0_6_54303)
  );
  LocalMux t4696 (
    .I(seg_11_15_sp4_v_b_17_42915),
    .O(seg_11_15_local_g0_1_46882)
  );
  Span4Mux_v3 t4697 (
    .I(seg_11_12_sp4_h_r_10_46608),
    .O(seg_11_15_sp4_v_b_17_42915)
  );
  LocalMux t4698 (
    .I(seg_13_14_sp4_r_v_b_7_54163),
    .O(seg_13_14_local_g1_7_54435)
  );
  LocalMux t4699 (
    .I(seg_13_13_lutff_0_out_50425),
    .O(seg_13_13_local_g2_0_54313)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t47 (
    .carryinitin(),
    .carryinitout(t46)
  );
  CascadeMux t470 (
    .I(net_34439),
    .O(net_34439_cascademuxed)
  );
  LocalMux t4700 (
    .I(seg_13_13_lutff_2_out_50427),
    .O(seg_13_13_local_g3_2_54323)
  );
  LocalMux t4701 (
    .I(seg_13_13_lutff_3_out_50428),
    .O(seg_13_13_local_g2_3_54316)
  );
  LocalMux t4702 (
    .I(seg_13_13_lutff_5_out_50430),
    .O(seg_13_13_local_g3_5_54326)
  );
  LocalMux t4703 (
    .I(seg_13_18_sp4_r_v_b_18_54778),
    .O(seg_13_18_local_g3_2_54938)
  );
  Span4Mux_v3 t4704 (
    .I(seg_14_15_sp4_v_b_7_54286),
    .O(seg_13_18_sp4_r_v_b_18_54778)
  );
  LocalMux t4705 (
    .I(seg_13_18_sp4_r_v_b_24_54896),
    .O(seg_13_18_local_g0_0_54912)
  );
  Span4Mux_v2 t4706 (
    .I(seg_14_16_sp4_v_b_4_54408),
    .O(seg_13_18_sp4_r_v_b_24_54896)
  );
  LocalMux t4707 (
    .I(seg_13_19_sp4_v_b_1_50941),
    .O(seg_13_19_local_g1_1_55044)
  );
  Span4Mux_v4 t4708 (
    .I(seg_13_15_sp4_v_b_10_50460),
    .O(seg_13_19_sp4_v_b_1_50941)
  );
  LocalMux t4709 (
    .I(seg_13_18_sp4_v_b_29_51068),
    .O(seg_13_18_local_g3_5_54941)
  );
  Span4Mux_v2 t4710 (
    .I(seg_13_16_sp4_v_b_9_50580),
    .O(seg_13_18_sp4_v_b_29_51068)
  );
  LocalMux t4711 (
    .I(seg_12_14_neigh_op_rgt_1_50549),
    .O(seg_12_14_local_g2_1_50606)
  );
  LocalMux t4712 (
    .I(seg_13_15_neigh_op_bot_1_50549),
    .O(seg_13_15_local_g1_1_54552)
  );
  LocalMux t4713 (
    .I(seg_14_14_neigh_op_lft_1_50549),
    .O(seg_14_14_local_g0_1_58251)
  );
  LocalMux t4714 (
    .I(seg_12_15_neigh_op_bnr_2_50550),
    .O(seg_12_15_local_g0_2_50714)
  );
  LocalMux t4715 (
    .I(seg_13_18_sp12_v_b_2_53651),
    .O(seg_13_18_local_g2_2_54930)
  );
  LocalMux t4716 (
    .I(seg_13_18_sp12_v_b_6_53897),
    .O(seg_13_18_local_g3_6_54942)
  );
  LocalMux t4717 (
    .I(seg_16_16_sp4_v_b_31_62315),
    .O(seg_16_16_local_g3_7_66188)
  );
  Span4Mux_v2 t4718 (
    .I(seg_16_14_sp4_h_l_42_50692),
    .O(seg_16_16_sp4_v_b_31_62315)
  );
  LocalMux t4719 (
    .I(seg_16_17_sp4_v_b_18_62315),
    .O(seg_16_17_local_g0_2_66282)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t472 (
    .carryinitin(),
    .carryinitout(t471)
  );
  Span4Mux_v3 t4720 (
    .I(seg_16_14_sp4_h_l_42_50692),
    .O(seg_16_17_sp4_v_b_18_62315)
  );
  LocalMux t4721 (
    .I(seg_17_14_sp4_h_r_14_66010),
    .O(seg_17_14_local_g0_6_69748)
  );
  Span4Mux_h1 t4722 (
    .I(seg_16_14_sp4_h_l_42_50692),
    .O(seg_17_14_sp4_h_r_14_66010)
  );
  LocalMux t4723 (
    .I(seg_20_12_sp4_v_b_25_76909),
    .O(seg_20_12_local_g3_1_80383)
  );
  Span4Mux_v2 t4724 (
    .I(seg_20_14_sp4_h_l_42_66014),
    .O(seg_20_12_sp4_v_b_25_76909)
  );
  Span4Mux_h4 t4725 (
    .I(seg_16_14_sp4_h_l_42_50692),
    .O(seg_20_14_sp4_h_l_42_66014)
  );
  LocalMux t4726 (
    .I(seg_16_17_sp4_r_v_b_15_66143),
    .O(seg_16_17_local_g2_7_66303)
  );
  Span4Mux_v3 t4727 (
    .I(seg_17_14_sp4_h_l_39_54518),
    .O(seg_16_17_sp4_r_v_b_15_66143)
  );
  LocalMux t4728 (
    .I(seg_17_14_sp4_h_r_5_69843),
    .O(seg_17_14_local_g0_5_69747)
  );
  Span4Mux_h0 t4729 (
    .I(seg_17_14_sp4_h_l_39_54518),
    .O(seg_17_14_sp4_h_r_5_69843)
  );
  CascadeMux t473 (
    .I(net_34562),
    .O(net_34562_cascademuxed)
  );
  LocalMux t4730 (
    .I(seg_17_17_sp4_v_b_15_66143),
    .O(seg_17_17_local_g0_7_70118)
  );
  Span4Mux_v3 t4731 (
    .I(seg_17_14_sp4_h_l_39_54518),
    .O(seg_17_17_sp4_v_b_15_66143)
  );
  LocalMux t4732 (
    .I(seg_11_18_sp4_v_b_10_43167),
    .O(seg_11_18_local_g1_2_47260)
  );
  Span4Mux_v4 t4733 (
    .I(seg_11_14_sp4_h_r_4_46858),
    .O(seg_11_18_sp4_v_b_10_43167)
  );
  LocalMux t4734 (
    .I(seg_10_18_sp4_r_v_b_4_43161),
    .O(seg_10_18_local_g1_4_43431)
  );
  Span4Mux_v4 t4735 (
    .I(seg_11_14_sp4_h_r_10_46854),
    .O(seg_10_18_sp4_r_v_b_4_43161)
  );
  LocalMux t4736 (
    .I(seg_11_12_sp4_v_b_34_42675),
    .O(seg_11_12_local_g3_2_46538)
  );
  Span4Mux_v2 t4737 (
    .I(seg_11_14_sp4_h_r_10_46854),
    .O(seg_11_12_sp4_v_b_34_42675)
  );
  LocalMux t4738 (
    .I(seg_13_18_sp4_r_v_b_5_54653),
    .O(seg_13_18_local_g1_5_54925)
  );
  Span4Mux_v4 t4739 (
    .I(seg_14_14_sp4_h_l_40_43028),
    .O(seg_13_18_sp4_r_v_b_5_54653)
  );
  CascadeMux t474 (
    .I(net_34568),
    .O(net_34568_cascademuxed)
  );
  LocalMux t4740 (
    .I(seg_13_8_sp4_r_v_b_35_53675),
    .O(seg_13_8_local_g0_0_53682)
  );
  Span4Mux_v2 t4741 (
    .I(seg_14_10_sp4_v_t_38_54159),
    .O(seg_13_8_sp4_r_v_b_35_53675)
  );
  LocalMux t4742 (
    .I(seg_14_18_sp4_v_b_3_54651),
    .O(seg_14_18_local_g1_3_58753)
  );
  Span4Mux_v4 t4743 (
    .I(seg_14_14_sp4_v_b_3_54159),
    .O(seg_14_18_sp4_v_b_3_54651)
  );
  LocalMux t4744 (
    .I(seg_15_10_sp4_h_r_14_57857),
    .O(seg_15_10_local_g0_6_61594)
  );
  Span4Mux_h1 t4745 (
    .I(seg_14_10_sp4_v_t_38_54159),
    .O(seg_15_10_sp4_h_r_14_57857)
  );
  LocalMux t4746 (
    .I(seg_11_16_sp4_h_r_22_43270),
    .O(seg_11_16_local_g1_6_47018)
  );
  Span4Mux_h3 t4747 (
    .I(seg_14_16_sp4_v_b_11_54413),
    .O(seg_11_16_sp4_h_r_22_43270)
  );
  LocalMux t4748 (
    .I(seg_14_18_sp4_v_b_26_54898),
    .O(seg_14_18_local_g3_2_58768)
  );
  Span4Mux_v2 t4749 (
    .I(seg_14_16_sp4_v_b_11_54413),
    .O(seg_14_18_sp4_v_b_26_54898)
  );
  CascadeMux t475 (
    .I(net_34574),
    .O(net_34574_cascademuxed)
  );
  LocalMux t4750 (
    .I(seg_13_18_sp4_v_b_8_50827),
    .O(seg_13_18_local_g1_0_54920)
  );
  Span4Mux_v4 t4751 (
    .I(seg_13_14_sp4_v_b_0_50327),
    .O(seg_13_18_sp4_v_b_8_50827)
  );
  LocalMux t4752 (
    .I(seg_13_18_sp4_v_b_43_51194),
    .O(seg_13_18_local_g2_3_54931)
  );
  Span4Mux_v1 t4753 (
    .I(seg_13_17_sp4_v_b_3_50697),
    .O(seg_13_18_sp4_v_b_43_51194)
  );
  LocalMux t4754 (
    .I(seg_13_16_neigh_op_bot_1_50672),
    .O(seg_13_16_local_g0_1_54667)
  );
  LocalMux t4755 (
    .I(seg_13_16_neigh_op_bot_2_50673),
    .O(seg_13_16_local_g1_2_54676)
  );
  GlobalMux t4756 (
    .I(seg_13_31_local_g1_0_56532_i3),
    .O(seg_10_18_glb_netwk_1_6)
  );
  gio2CtrlBuf t4757 (
    .I(seg_13_31_local_g1_0_56532_i2),
    .O(seg_13_31_local_g1_0_56532_i3)
  );
  ICE_GB t4758 (
    .GLOBALBUFFEROUTPUT(seg_13_31_local_g1_0_56532_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_13_31_local_g1_0_56532_i1)
  );
  IoInMux t4759 (
    .I(seg_13_31_local_g1_0_56532),
    .O(seg_13_31_local_g1_0_56532_i1)
  );
  CascadeMux t476 (
    .I(net_34580),
    .O(net_34580_cascademuxed)
  );
  LocalMux t4760 (
    .I(seg_13_31_span12_vert_8_55620),
    .O(seg_13_31_local_g1_0_56532)
  );
  Span12Mux_v8 t4761 (
    .I(seg_13_23_sp12_v_b_0_54144),
    .O(seg_13_31_span12_vert_8_55620)
  );
  LocalMux t4762 (
    .I(seg_13_18_sp4_r_v_b_4_54654),
    .O(seg_13_18_local_g1_4_54924)
  );
  LocalMux t4763 (
    .I(seg_13_18_sp4_r_v_b_6_54656),
    .O(seg_13_18_local_g1_6_54926)
  );
  LocalMux t4764 (
    .I(seg_13_18_sp4_r_v_b_8_54658),
    .O(seg_13_18_local_g2_0_54928)
  );
  LocalMux t4765 (
    .I(seg_12_13_sp4_r_v_b_42_50578),
    .O(seg_12_13_local_g3_2_50492)
  );
  LocalMux t4766 (
    .I(seg_13_18_sp4_v_b_11_50828),
    .O(seg_13_18_local_g0_3_54915)
  );
  LocalMux t4767 (
    .I(seg_13_15_neigh_op_top_1_50795),
    .O(seg_13_15_local_g0_1_54544)
  );
  LocalMux t4768 (
    .I(seg_13_16_lutff_2_out_50796),
    .O(seg_13_16_local_g0_2_54668)
  );
  LocalMux t4769 (
    .I(seg_12_15_neigh_op_tnr_3_50797),
    .O(seg_12_15_local_g2_3_50731)
  );
  CascadeMux t477 (
    .I(net_34586),
    .O(net_34586_cascademuxed)
  );
  LocalMux t4770 (
    .I(seg_13_15_neigh_op_top_3_50797),
    .O(seg_13_15_local_g0_3_54546)
  );
  LocalMux t4771 (
    .I(seg_13_16_lutff_3_out_50797),
    .O(seg_13_16_local_g2_3_54685)
  );
  LocalMux t4772 (
    .I(seg_13_17_neigh_op_bot_3_50797),
    .O(seg_13_17_local_g1_3_54800)
  );
  LocalMux t4773 (
    .I(seg_13_16_lutff_4_out_50798),
    .O(seg_13_16_local_g3_4_54694)
  );
  LocalMux t4774 (
    .I(seg_13_16_lutff_5_out_50799),
    .O(seg_13_16_local_g3_5_54695)
  );
  LocalMux t4775 (
    .I(seg_13_15_neigh_op_top_6_50800),
    .O(seg_13_15_local_g0_6_54549)
  );
  LocalMux t4776 (
    .I(seg_12_16_neigh_op_rgt_7_50801),
    .O(seg_12_16_local_g2_7_50858)
  );
  LocalMux t4777 (
    .I(seg_13_16_lutff_7_out_50801),
    .O(seg_13_16_local_g0_7_54673)
  );
  LocalMux t4778 (
    .I(seg_11_18_sp4_r_v_b_26_47236),
    .O(seg_11_18_local_g0_2_47252)
  );
  Span4Mux_v2 t4779 (
    .I(seg_12_16_sp4_v_b_11_46751),
    .O(seg_11_18_sp4_r_v_b_26_47236)
  );
  CascadeMux t478 (
    .I(net_34592),
    .O(net_34592_cascademuxed)
  );
  Span4Mux_v0 t4780 (
    .I(seg_12_16_sp4_h_r_11_50932),
    .O(seg_12_16_sp4_v_b_11_46751)
  );
  LocalMux t4781 (
    .I(seg_16_12_sp4_h_r_10_65761),
    .O(seg_16_12_local_g0_2_65667)
  );
  Span4Mux_h0 t4782 (
    .I(seg_16_12_sp4_v_t_40_62067),
    .O(seg_16_12_sp4_h_r_10_65761)
  );
  Span4Mux_v4 t4783 (
    .I(seg_16_16_sp4_h_l_46_50932),
    .O(seg_16_12_sp4_v_t_40_62067)
  );
  LocalMux t4784 (
    .I(seg_9_18_sp4_r_v_b_27_39573),
    .O(seg_9_18_local_g1_3_39599)
  );
  Span4Mux_v2 t4785 (
    .I(seg_10_16_sp4_h_r_3_43272),
    .O(seg_9_18_sp4_r_v_b_27_39573)
  );
  LocalMux t4786 (
    .I(seg_13_18_sp4_r_v_b_27_54897),
    .O(seg_13_18_local_g1_3_54923)
  );
  Span4Mux_v2 t4787 (
    .I(seg_14_16_sp4_h_l_38_43272),
    .O(seg_13_18_sp4_r_v_b_27_54897)
  );
  LocalMux t4788 (
    .I(seg_8_15_sp4_h_r_26_28139),
    .O(seg_8_15_local_g2_2_35406)
  );
  Span4Mux_h2 t4789 (
    .I(seg_10_15_sp4_h_r_2_43148),
    .O(seg_8_15_sp4_h_r_26_28139)
  );
  CascadeMux t479 (
    .I(net_34598),
    .O(net_34598_cascademuxed)
  );
  Span4Mux_h4 t4790 (
    .I(seg_14_15_sp4_v_t_39_54775),
    .O(seg_10_15_sp4_h_r_2_43148)
  );
  LocalMux t4791 (
    .I(seg_17_8_sp4_h_r_42_57615),
    .O(seg_17_8_local_g2_2_69022)
  );
  Span4Mux_h3 t4792 (
    .I(seg_14_8_sp4_v_t_42_53917),
    .O(seg_17_8_sp4_h_r_42_57615)
  );
  Span4Mux_v4 t4793 (
    .I(seg_14_12_sp4_v_t_42_54409),
    .O(seg_14_8_sp4_v_t_42_53917)
  );
  LocalMux t4794 (
    .I(seg_14_13_sp4_v_b_44_54411),
    .O(seg_14_13_local_g3_4_58155)
  );
  LocalMux t4795 (
    .I(seg_14_14_sp4_v_b_33_54411),
    .O(seg_14_14_local_g3_1_58275)
  );
  LocalMux t4796 (
    .I(seg_13_19_sp4_v_b_3_50943),
    .O(seg_13_19_local_g1_3_55046)
  );
  LocalMux t4797 (
    .I(seg_13_17_lutff_1_out_50918),
    .O(seg_13_17_local_g0_1_54790)
  );
  LocalMux t4798 (
    .I(seg_13_16_neigh_op_top_3_50920),
    .O(seg_13_16_local_g0_3_54669)
  );
  LocalMux t4799 (
    .I(seg_13_16_neigh_op_top_3_50920),
    .O(seg_13_16_local_g1_3_54677)
  );
  CascadeMux t48 (
    .I(net_8854),
    .O(net_8854_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t480 (
    .carryinitin(net_38432),
    .carryinitout(net_38476)
  );
  LocalMux t4800 (
    .I(seg_13_17_lutff_3_out_50920),
    .O(seg_13_17_local_g3_3_54816)
  );
  LocalMux t4801 (
    .I(seg_13_16_neigh_op_top_4_50921),
    .O(seg_13_16_local_g1_4_54678)
  );
  LocalMux t4802 (
    .I(seg_13_17_lutff_4_out_50921),
    .O(seg_13_17_local_g0_4_54793)
  );
  LocalMux t4803 (
    .I(seg_12_16_neigh_op_tnr_5_50922),
    .O(seg_12_16_local_g3_5_50864)
  );
  LocalMux t4804 (
    .I(seg_13_16_neigh_op_top_5_50922),
    .O(seg_13_16_local_g1_5_54679)
  );
  LocalMux t4805 (
    .I(seg_12_16_neigh_op_tnr_7_50924),
    .O(seg_12_16_local_g3_7_50866)
  );
  LocalMux t4806 (
    .I(seg_13_17_lutff_7_out_50924),
    .O(seg_13_17_local_g0_7_54796)
  );
  LocalMux t4807 (
    .I(seg_13_18_neigh_op_bot_7_50924),
    .O(seg_13_18_local_g1_7_54927)
  );
  LocalMux t4808 (
    .I(seg_16_12_sp4_v_b_13_61695),
    .O(seg_16_12_local_g1_5_65678)
  );
  Span4Mux_v1 t4809 (
    .I(seg_16_13_sp4_v_t_44_62194),
    .O(seg_16_12_sp4_v_b_13_61695)
  );
  CascadeMux t481 (
    .I(net_34691),
    .O(net_34691_cascademuxed)
  );
  Span4Mux_v4 t4810 (
    .I(seg_16_17_sp4_h_l_38_51057),
    .O(seg_16_13_sp4_v_t_44_62194)
  );
  LocalMux t4811 (
    .I(seg_9_13_sp4_h_r_30_31413),
    .O(seg_9_13_local_g3_6_39003)
  );
  Span4Mux_h2 t4812 (
    .I(seg_11_13_sp4_v_t_43_43040),
    .O(seg_9_13_sp4_h_r_30_31413)
  );
  Span4Mux_v4 t4813 (
    .I(seg_11_17_sp4_h_r_6_47229),
    .O(seg_11_13_sp4_v_t_43_43040)
  );
  LocalMux t4814 (
    .I(seg_10_11_sp4_r_v_b_26_42544),
    .O(seg_10_11_local_g0_2_42560)
  );
  Span4Mux_v2 t4815 (
    .I(seg_11_13_sp4_v_t_43_43040),
    .O(seg_10_11_sp4_r_v_b_26_42544)
  );
  LocalMux t4816 (
    .I(seg_11_12_sp4_v_b_15_42544),
    .O(seg_11_12_local_g1_7_46527)
  );
  Span4Mux_v1 t4817 (
    .I(seg_11_13_sp4_v_t_43_43040),
    .O(seg_11_12_sp4_v_b_15_42544)
  );
  LocalMux t4818 (
    .I(seg_9_14_sp4_r_v_b_46_39212),
    .O(seg_9_14_local_g3_6_39126)
  );
  Span4Mux_v3 t4819 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_9_14_sp4_r_v_b_46_39212)
  );
  CascadeMux t482 (
    .I(net_34709),
    .O(net_34709_cascademuxed)
  );
  LocalMux t4820 (
    .I(seg_9_17_sp4_r_v_b_11_39212),
    .O(seg_9_17_local_g2_3_39484)
  );
  Span4Mux_v1 t4821 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_9_17_sp4_r_v_b_11_39212)
  );
  LocalMux t4822 (
    .I(seg_9_18_sp4_r_v_b_40_39698),
    .O(seg_9_18_local_g3_0_39612)
  );
  Span4Mux_v1 t4823 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_9_18_sp4_r_v_b_40_39698)
  );
  LocalMux t4824 (
    .I(seg_10_15_sp4_v_b_35_39212),
    .O(seg_10_15_local_g3_3_43077)
  );
  Span4Mux_v2 t4825 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_10_15_sp4_v_b_35_39212)
  );
  LocalMux t4826 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_10_17_local_g0_3_43299)
  );
  LocalMux t4827 (
    .I(seg_11_13_sp4_h_r_17_42904),
    .O(seg_11_13_local_g0_1_46636)
  );
  Span4Mux_h1 t4828 (
    .I(seg_10_13_sp4_v_t_46_39212),
    .O(seg_11_13_sp4_h_r_17_42904)
  );
  Span4Mux_v4 t4829 (
    .I(seg_10_17_sp4_h_r_11_43393),
    .O(seg_10_13_sp4_v_t_46_39212)
  );
  CascadeMux t483 (
    .I(net_34820),
    .O(net_34820_cascademuxed)
  );
  LocalMux t4830 (
    .I(seg_11_17_sp4_h_r_22_43393),
    .O(seg_11_17_local_g1_6_47141)
  );
  LocalMux t4831 (
    .I(seg_11_18_sp4_h_r_15_43517),
    .O(seg_11_18_local_g0_7_47257)
  );
  Span4Mux_h3 t4832 (
    .I(seg_14_18_sp4_v_b_2_54652),
    .O(seg_11_18_sp4_h_r_15_43517)
  );
  LocalMux t4833 (
    .I(seg_11_18_sp4_h_r_15_43517),
    .O(seg_11_18_local_g1_7_47265)
  );
  LocalMux t4834 (
    .I(seg_14_8_sp4_v_b_29_53669),
    .O(seg_14_8_local_g3_5_57541)
  );
  Span4Mux_v2 t4835 (
    .I(seg_14_10_sp4_v_t_39_54160),
    .O(seg_14_8_sp4_v_b_29_53669)
  );
  Span4Mux_v4 t4836 (
    .I(seg_14_14_sp4_v_t_39_54652),
    .O(seg_14_10_sp4_v_t_39_54160)
  );
  LocalMux t4837 (
    .I(seg_14_9_sp4_v_b_16_53669),
    .O(seg_14_9_local_g1_0_57643)
  );
  Span4Mux_v1 t4838 (
    .I(seg_14_10_sp4_v_t_39_54160),
    .O(seg_14_9_sp4_v_b_16_53669)
  );
  LocalMux t4839 (
    .I(seg_9_18_sp4_h_r_8_39692),
    .O(seg_9_18_local_g0_0_39588)
  );
  CascadeMux t484 (
    .I(net_34937),
    .O(net_34937_cascademuxed)
  );
  Span4Mux_h4 t4840 (
    .I(seg_13_18_sp4_v_b_3_50820),
    .O(seg_9_18_sp4_h_r_8_39692)
  );
  LocalMux t4841 (
    .I(seg_12_12_sp4_r_v_b_35_50336),
    .O(seg_12_12_local_g2_3_50362)
  );
  Span4Mux_v2 t4842 (
    .I(seg_13_14_sp4_v_t_38_50820),
    .O(seg_12_12_sp4_r_v_b_35_50336)
  );
  LocalMux t4843 (
    .I(seg_13_8_sp4_v_b_35_49844),
    .O(seg_13_8_local_g2_3_53701)
  );
  Span4Mux_v2 t4844 (
    .I(seg_13_10_sp4_v_t_46_50336),
    .O(seg_13_8_sp4_v_b_35_49844)
  );
  Span4Mux_v4 t4845 (
    .I(seg_13_14_sp4_v_t_38_50820),
    .O(seg_13_10_sp4_v_t_46_50336)
  );
  LocalMux t4846 (
    .I(seg_13_10_sp4_h_r_4_54028),
    .O(seg_13_10_local_g1_4_53940)
  );
  Span4Mux_h0 t4847 (
    .I(seg_13_10_sp4_v_t_46_50336),
    .O(seg_13_10_sp4_h_r_4_54028)
  );
  LocalMux t4848 (
    .I(seg_13_11_sp4_v_b_46_50336),
    .O(seg_13_11_local_g2_6_54073)
  );
  Span4Mux_v3 t4849 (
    .I(seg_13_14_sp4_v_t_38_50820),
    .O(seg_13_11_sp4_v_b_46_50336)
  );
  CascadeMux t485 (
    .I(net_35054),
    .O(net_35054_cascademuxed)
  );
  LocalMux t4850 (
    .I(seg_13_13_sp4_v_b_22_50336),
    .O(seg_13_13_local_g1_6_54311)
  );
  Span4Mux_v1 t4851 (
    .I(seg_13_14_sp4_v_t_38_50820),
    .O(seg_13_13_sp4_v_b_22_50336)
  );
  LocalMux t4852 (
    .I(seg_13_14_sp4_h_r_8_54524),
    .O(seg_13_14_local_g1_0_54428)
  );
  Span4Mux_h0 t4853 (
    .I(seg_13_14_sp4_v_t_38_50820),
    .O(seg_13_14_sp4_h_r_8_54524)
  );
  LocalMux t4854 (
    .I(seg_17_8_sp4_v_b_28_65161),
    .O(seg_17_8_local_g2_4_69024)
  );
  Span4Mux_v2 t4855 (
    .I(seg_17_10_sp4_h_l_41_54028),
    .O(seg_17_8_sp4_v_b_28_65161)
  );
  Span4Mux_h4 t4856 (
    .I(seg_13_10_sp4_v_t_46_50336),
    .O(seg_17_10_sp4_h_l_41_54028)
  );
  LocalMux t4857 (
    .I(seg_17_8_sp4_v_b_28_65161),
    .O(seg_17_8_local_g3_4_69032)
  );
  LocalMux t4858 (
    .I(seg_8_15_sp4_r_v_b_11_35135),
    .O(seg_8_15_local_g2_3_35407)
  );
  Span4Mux_v1 t4859 (
    .I(seg_9_15_sp4_h_r_6_39321),
    .O(seg_8_15_sp4_r_v_b_11_35135)
  );
  CascadeMux t486 (
    .I(net_35066),
    .O(net_35066_cascademuxed)
  );
  Span4Mux_h4 t4860 (
    .I(seg_13_15_sp4_v_t_43_50948),
    .O(seg_9_15_sp4_h_r_6_39321)
  );
  LocalMux t4861 (
    .I(seg_9_15_sp4_h_r_6_39321),
    .O(seg_9_15_local_g1_6_39233)
  );
  LocalMux t4862 (
    .I(seg_11_11_sp4_h_r_24_38821),
    .O(seg_11_11_local_g2_0_46405)
  );
  Span4Mux_h2 t4863 (
    .I(seg_13_11_sp4_v_t_43_50456),
    .O(seg_11_11_sp4_h_r_24_38821)
  );
  Span4Mux_v4 t4864 (
    .I(seg_13_15_sp4_v_t_43_50948),
    .O(seg_13_11_sp4_v_t_43_50456)
  );
  LocalMux t4865 (
    .I(seg_11_15_sp4_h_r_30_39321),
    .O(seg_11_15_local_g3_6_46911)
  );
  Span4Mux_h2 t4866 (
    .I(seg_13_15_sp4_v_t_43_50948),
    .O(seg_11_15_sp4_h_r_30_39321)
  );
  LocalMux t4867 (
    .I(seg_13_19_sp4_v_b_6_50948),
    .O(seg_13_19_local_g1_6_55049)
  );
  LocalMux t4868 (
    .I(seg_14_18_neigh_op_lft_1_51041),
    .O(seg_14_18_local_g0_1_58743)
  );
  LocalMux t4869 (
    .I(seg_14_18_neigh_op_lft_2_51042),
    .O(seg_14_18_local_g1_2_58752)
  );
  CascadeMux t487 (
    .I(net_35078),
    .O(net_35078_cascademuxed)
  );
  LocalMux t4870 (
    .I(seg_14_18_neigh_op_lft_6_51046),
    .O(seg_14_18_local_g0_6_58748)
  );
  LocalMux t4871 (
    .I(seg_12_14_sp4_h_r_1_50684),
    .O(seg_12_14_local_g1_1_50598)
  );
  Span4Mux_h0 t4872 (
    .I(seg_12_14_sp4_v_t_45_46996),
    .O(seg_12_14_sp4_h_r_1_50684)
  );
  Span4Mux_v4 t4873 (
    .I(seg_12_18_sp4_h_r_3_51180),
    .O(seg_12_14_sp4_v_t_45_46996)
  );
  LocalMux t4874 (
    .I(seg_10_18_sp4_h_r_3_43518),
    .O(seg_10_18_local_g0_3_43422)
  );
  LocalMux t4875 (
    .I(seg_11_16_sp4_h_r_26_39440),
    .O(seg_11_16_local_g2_2_47022)
  );
  Span4Mux_h2 t4876 (
    .I(seg_13_16_sp4_v_t_39_51067),
    .O(seg_11_16_sp4_h_r_26_39440)
  );
  LocalMux t4877 (
    .I(seg_11_12_sp4_h_r_28_38950),
    .O(seg_11_12_local_g3_4_46540)
  );
  Span4Mux_h2 t4878 (
    .I(seg_13_12_sp4_v_t_41_50577),
    .O(seg_11_12_sp4_h_r_28_38950)
  );
  Span4Mux_v4 t4879 (
    .I(seg_13_16_sp4_v_t_45_51073),
    .O(seg_13_12_sp4_v_t_41_50577)
  );
  CascadeMux t488 (
    .I(net_35189),
    .O(net_35189_cascademuxed)
  );
  LocalMux t4880 (
    .I(seg_11_16_sp4_h_r_27_39441),
    .O(seg_11_16_local_g3_3_47031)
  );
  Span4Mux_h2 t4881 (
    .I(seg_13_16_sp4_v_t_38_51066),
    .O(seg_11_16_sp4_h_r_27_39441)
  );
  GlobalMux t4882 (
    .I(seg_19_0_local_g1_0_75715_i3),
    .O(seg_3_8_glb_netwk_7_12)
  );
  gio2CtrlBuf t4883 (
    .I(seg_19_0_local_g1_0_75715_i2),
    .O(seg_19_0_local_g1_0_75715_i3)
  );
  ICE_GB t4884 (
    .GLOBALBUFFEROUTPUT(seg_19_0_local_g1_0_75715_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_19_0_local_g1_0_75715_i1)
  );
  IoInMux t4885 (
    .I(seg_19_0_local_g1_0_75715),
    .O(seg_19_0_local_g1_0_75715_i1)
  );
  LocalMux t4886 (
    .I(seg_19_0_span4_vert_0_72044),
    .O(seg_19_0_local_g1_0_75715)
  );
  Span4Mux_v1 t4887 (
    .I(seg_19_1_sp4_h_l_37_60539),
    .O(seg_19_0_span4_vert_0_72044)
  );
  Span4Mux_h4 t4888 (
    .I(seg_15_1_sp4_h_l_44_45228),
    .O(seg_19_1_sp4_h_l_37_60539)
  );
  LocalMux t4889 (
    .I(seg_14_2_lutff_0_out_52867),
    .O(seg_14_2_local_g0_0_56774)
  );
  CascadeMux t489 (
    .I(net_35207),
    .O(net_35207_cascademuxed)
  );
  LocalMux t4890 (
    .I(seg_14_2_lutff_2_out_52869),
    .O(seg_14_2_local_g0_2_56776)
  );
  LocalMux t4891 (
    .I(seg_14_2_lutff_6_out_52873),
    .O(seg_14_2_local_g1_6_56788)
  );
  LocalMux t4892 (
    .I(seg_14_4_sp4_r_v_b_15_56883),
    .O(seg_14_4_local_g2_7_57043)
  );
  LocalMux t4893 (
    .I(seg_14_4_neigh_op_bot_6_53032),
    .O(seg_14_4_local_g0_6_57026)
  );
  LocalMux t4894 (
    .I(seg_14_4_neigh_op_bot_7_53033),
    .O(seg_14_4_local_g1_7_57035)
  );
  LocalMux t4895 (
    .I(seg_14_5_neigh_op_bot_0_53149),
    .O(seg_14_5_local_g0_0_57143)
  );
  LocalMux t4896 (
    .I(seg_13_3_neigh_op_tnr_2_53151),
    .O(seg_13_3_local_g3_2_53093)
  );
  LocalMux t4897 (
    .I(seg_15_4_neigh_op_lft_2_53151),
    .O(seg_15_4_local_g0_2_60852)
  );
  LocalMux t4898 (
    .I(seg_15_5_neigh_op_bnl_2_53151),
    .O(seg_15_5_local_g2_2_60991)
  );
  LocalMux t4899 (
    .I(seg_14_5_neigh_op_bot_3_53152),
    .O(seg_14_5_local_g0_3_57146)
  );
  CascadeMux t49 (
    .I(net_8866),
    .O(net_8866_cascademuxed)
  );
  CascadeMux t490 (
    .I(net_35336),
    .O(net_35336_cascademuxed)
  );
  LocalMux t4900 (
    .I(seg_14_5_neigh_op_bot_5_53154),
    .O(seg_14_5_local_g1_5_57156)
  );
  LocalMux t4901 (
    .I(seg_12_10_sp4_r_v_b_24_50081),
    .O(seg_12_10_local_g0_0_50097)
  );
  Span4Mux_v2 t4902 (
    .I(seg_13_8_sp4_v_b_9_49596),
    .O(seg_12_10_sp4_r_v_b_24_50081)
  );
  Span4Mux_v4 t4903 (
    .I(seg_13_4_sp4_h_r_9_53295),
    .O(seg_13_8_sp4_v_b_9_49596)
  );
  LocalMux t4904 (
    .I(seg_16_10_sp4_r_v_b_24_65403),
    .O(seg_16_10_local_g1_0_65427)
  );
  Span4Mux_v2 t4905 (
    .I(seg_17_8_sp4_v_b_9_64918),
    .O(seg_16_10_sp4_r_v_b_24_65403)
  );
  Span4Mux_v4 t4906 (
    .I(seg_17_4_sp4_h_l_44_53295),
    .O(seg_17_8_sp4_v_b_9_64918)
  );
  LocalMux t4907 (
    .I(seg_12_4_sp4_h_r_6_49461),
    .O(seg_12_4_local_g1_6_49373)
  );
  LocalMux t4908 (
    .I(seg_11_2_sp4_v_b_30_41436),
    .O(seg_11_2_local_g3_6_45312)
  );
  Span4Mux_v2 t4909 (
    .I(seg_11_4_sp4_h_r_1_45623),
    .O(seg_11_2_sp4_v_b_30_41436)
  );
  CascadeMux t491 (
    .I(net_35423),
    .O(net_35423_cascademuxed)
  );
  LocalMux t4910 (
    .I(seg_12_13_sp4_h_r_18_46738),
    .O(seg_12_13_local_g1_2_50476)
  );
  Span4Mux_h3 t4911 (
    .I(seg_15_13_sp4_v_b_2_57867),
    .O(seg_12_13_sp4_h_r_18_46738)
  );
  Span4Mux_v4 t4912 (
    .I(seg_15_9_sp4_v_b_11_57382),
    .O(seg_15_13_sp4_v_b_2_57867)
  );
  Span4Mux_v4 t4913 (
    .I(seg_15_5_sp4_v_b_8_56889),
    .O(seg_15_9_sp4_v_b_11_57382)
  );
  LocalMux t4914 (
    .I(seg_14_6_sp4_r_v_b_1_57003),
    .O(seg_14_6_local_g1_1_57275)
  );
  LocalMux t4915 (
    .I(seg_14_6_sp4_r_v_b_21_57135),
    .O(seg_14_6_local_g3_5_57295)
  );
  LocalMux t4916 (
    .I(seg_14_6_sp4_v_b_12_53296),
    .O(seg_14_6_local_g0_4_57270)
  );
  LocalMux t4917 (
    .I(seg_14_10_sp4_v_b_17_53793),
    .O(seg_14_10_local_g0_1_57759)
  );
  Span4Mux_v3 t4918 (
    .I(seg_14_7_sp4_v_b_1_53296),
    .O(seg_14_10_sp4_v_b_17_53793)
  );
  LocalMux t4919 (
    .I(seg_14_5_lutff_1_out_53273),
    .O(seg_14_5_local_g2_1_57160)
  );
  CascadeMux t492 (
    .I(net_35429),
    .O(net_35429_cascademuxed)
  );
  LocalMux t4920 (
    .I(seg_14_5_lutff_2_out_53274),
    .O(seg_14_5_local_g0_2_57145)
  );
  LocalMux t4921 (
    .I(seg_14_6_neigh_op_bot_3_53275),
    .O(seg_14_6_local_g0_3_57269)
  );
  LocalMux t4922 (
    .I(seg_15_6_neigh_op_bnl_4_53276),
    .O(seg_15_6_local_g3_4_61124)
  );
  LocalMux t4923 (
    .I(seg_15_6_neigh_op_bnl_5_53277),
    .O(seg_15_6_local_g3_5_61125)
  );
  LocalMux t4924 (
    .I(seg_14_5_lutff_6_out_53278),
    .O(seg_14_5_local_g3_6_57173)
  );
  LocalMux t4925 (
    .I(seg_14_6_neigh_op_bot_7_53279),
    .O(seg_14_6_local_g0_7_57273)
  );
  LocalMux t4926 (
    .I(seg_20_6_sp4_h_r_18_76396),
    .O(seg_20_6_local_g1_2_79630)
  );
  Span4Mux_h1 t4927 (
    .I(seg_19_6_sp4_h_l_41_61196),
    .O(seg_20_6_sp4_h_r_18_76396)
  );
  Span4Mux_h4 t4928 (
    .I(seg_15_6_sp4_v_b_4_57008),
    .O(seg_19_6_sp4_h_l_41_61196)
  );
  LocalMux t4929 (
    .I(seg_14_6_lutff_0_out_53395),
    .O(seg_14_6_local_g0_0_57266)
  );
  CascadeMux t493 (
    .I(net_35435),
    .O(net_35435_cascademuxed)
  );
  LocalMux t4930 (
    .I(seg_15_6_neigh_op_lft_3_53398),
    .O(seg_15_6_local_g0_3_61099)
  );
  LocalMux t4931 (
    .I(seg_14_7_neigh_op_bot_5_53400),
    .O(seg_14_7_local_g1_5_57402)
  );
  LocalMux t4932 (
    .I(seg_15_6_neigh_op_lft_7_53402),
    .O(seg_15_6_local_g1_7_61111)
  );
  LocalMux t4933 (
    .I(seg_25_7_sp4_v_b_39_95260),
    .O(seg_25_7_local_g2_7_99543)
  );
  Span4Mux_v1 t4934 (
    .I(seg_25_6_sp4_h_l_44_83556),
    .O(seg_25_7_sp4_v_b_39_95260)
  );
  Sp12to4 t4935 (
    .I(seg_22_6_sp12_h_r_16_57356),
    .O(seg_25_6_sp4_h_l_44_83556)
  );
  LocalMux t4936 (
    .I(seg_20_6_sp4_h_r_34_72685),
    .O(seg_20_6_local_g3_2_79646)
  );
  Span4Mux_h2 t4937 (
    .I(seg_18_6_sp4_h_l_39_57364),
    .O(seg_20_6_sp4_h_r_34_72685)
  );
  LocalMux t4938 (
    .I(seg_12_6_sp4_h_r_20_45879),
    .O(seg_12_6_local_g1_4_49617)
  );
  LocalMux t4939 (
    .I(seg_25_6_sp4_h_r_46_87379),
    .O(seg_25_6_local_g3_6_99400)
  );
  CascadeMux t494 (
    .I(net_35441),
    .O(net_35441_cascademuxed)
  );
  Span4Mux_h3 t4940 (
    .I(seg_22_6_sp4_h_l_46_72686),
    .O(seg_25_6_sp4_h_r_46_87379)
  );
  Span4Mux_h4 t4941 (
    .I(seg_18_6_sp4_h_l_45_57370),
    .O(seg_22_6_sp4_h_l_46_72686)
  );
  LocalMux t4942 (
    .I(seg_14_8_neigh_op_bot_1_53519),
    .O(seg_14_8_local_g1_1_57521)
  );
  LocalMux t4943 (
    .I(seg_14_8_neigh_op_bot_5_53523),
    .O(seg_14_8_local_g1_5_57525)
  );
  LocalMux t4944 (
    .I(seg_13_7_neigh_op_rgt_6_53524),
    .O(seg_13_7_local_g3_6_53589)
  );
  LocalMux t4945 (
    .I(seg_14_7_lutff_7_out_53525),
    .O(seg_14_7_local_g0_7_57396)
  );
  LocalMux t4946 (
    .I(seg_13_11_sp4_v_b_7_49963),
    .O(seg_13_11_local_g1_7_54066)
  );
  Span4Mux_v4 t4947 (
    .I(seg_13_7_sp4_h_r_1_53654),
    .O(seg_13_11_sp4_v_b_7_49963)
  );
  LocalMux t4948 (
    .I(seg_12_11_sp4_v_b_4_46131),
    .O(seg_12_11_local_g0_4_50224)
  );
  Span4Mux_v4 t4949 (
    .I(seg_12_7_sp4_h_r_4_49828),
    .O(seg_12_11_sp4_v_b_4_46131)
  );
  CascadeMux t495 (
    .I(net_35447),
    .O(net_35447_cascademuxed)
  );
  LocalMux t4950 (
    .I(seg_10_7_sp4_r_v_b_8_41812),
    .O(seg_10_7_local_g2_0_42082)
  );
  Span4Mux_v1 t4951 (
    .I(seg_11_7_sp4_h_r_3_45996),
    .O(seg_10_7_sp4_r_v_b_8_41812)
  );
  LocalMux t4952 (
    .I(seg_13_10_sp4_r_v_b_9_53673),
    .O(seg_13_10_local_g2_1_53945)
  );
  LocalMux t4953 (
    .I(seg_15_8_neigh_op_lft_5_53646),
    .O(seg_15_8_local_g1_5_61355)
  );
  LocalMux t4954 (
    .I(seg_11_8_sp4_h_r_21_42293),
    .O(seg_11_8_local_g0_5_46025)
  );
  Span4Mux_h3 t4955 (
    .I(seg_14_8_sp4_h_r_0_57606),
    .O(seg_11_8_sp4_h_r_21_42293)
  );
  LocalMux t4956 (
    .I(seg_17_8_sp4_h_r_1_69099),
    .O(seg_17_8_local_g0_1_69005)
  );
  Span4Mux_h0 t4957 (
    .I(seg_17_8_sp4_h_l_36_53777),
    .O(seg_17_8_sp4_h_r_1_69099)
  );
  LocalMux t4958 (
    .I(seg_11_8_sp4_h_r_16_42290),
    .O(seg_11_8_local_g1_0_46028)
  );
  Span4Mux_h3 t4959 (
    .I(seg_14_8_sp4_h_r_2_57610),
    .O(seg_11_8_sp4_h_r_16_42290)
  );
  CascadeMux t496 (
    .I(net_35459),
    .O(net_35459_cascademuxed)
  );
  LocalMux t4960 (
    .I(seg_12_18_sp4_r_v_b_25_51064),
    .O(seg_12_18_local_g0_1_51082)
  );
  Span4Mux_v2 t4961 (
    .I(seg_13_16_sp4_v_b_5_50576),
    .O(seg_12_18_sp4_r_v_b_25_51064)
  );
  Span4Mux_v4 t4962 (
    .I(seg_13_12_sp4_v_b_5_50084),
    .O(seg_13_16_sp4_v_b_5_50576)
  );
  Span4Mux_v4 t4963 (
    .I(seg_13_8_sp4_h_r_11_53779),
    .O(seg_13_12_sp4_v_b_5_50084)
  );
  LocalMux t4964 (
    .I(seg_11_15_sp4_v_b_20_42918),
    .O(seg_11_15_local_g0_4_46885)
  );
  Span4Mux_v3 t4965 (
    .I(seg_11_12_sp4_v_b_9_42426),
    .O(seg_11_15_sp4_v_b_20_42918)
  );
  Span4Mux_v4 t4966 (
    .I(seg_11_8_sp4_h_r_3_46119),
    .O(seg_11_12_sp4_v_b_9_42426)
  );
  LocalMux t4967 (
    .I(seg_11_8_sp4_h_r_5_46121),
    .O(seg_11_8_local_g1_5_46033)
  );
  LocalMux t4968 (
    .I(seg_10_11_sp4_r_v_b_22_42428),
    .O(seg_10_11_local_g3_6_42588)
  );
  Span4Mux_v3 t4969 (
    .I(seg_11_8_sp4_h_r_11_46117),
    .O(seg_10_11_sp4_r_v_b_22_42428)
  );
  CascadeMux t497 (
    .I(net_35465),
    .O(net_35465_cascademuxed)
  );
  LocalMux t4970 (
    .I(seg_11_10_sp4_v_b_35_42428),
    .O(seg_11_10_local_g2_3_46285)
  );
  Span4Mux_v2 t4971 (
    .I(seg_11_8_sp4_h_r_11_46117),
    .O(seg_11_10_sp4_v_b_35_42428)
  );
  LocalMux t4972 (
    .I(seg_11_14_sp4_v_b_21_42796),
    .O(seg_11_14_local_g1_5_46771)
  );
  Span4Mux_v3 t4973 (
    .I(seg_11_11_sp4_h_r_2_46487),
    .O(seg_11_14_sp4_v_b_21_42796)
  );
  Span4Mux_h4 t4974 (
    .I(seg_15_11_sp4_v_b_2_57621),
    .O(seg_11_11_sp4_h_r_2_46487)
  );
  LocalMux t4975 (
    .I(seg_12_11_sp4_h_r_23_46485),
    .O(seg_12_11_local_g0_7_50227)
  );
  Span4Mux_h3 t4976 (
    .I(seg_15_11_sp4_v_b_10_57629),
    .O(seg_12_11_sp4_h_r_23_46485)
  );
  LocalMux t4977 (
    .I(seg_9_12_sp4_r_v_b_15_38713),
    .O(seg_9_12_local_g2_7_38873)
  );
  Span4Mux_v3 t4978 (
    .I(seg_10_9_sp4_h_r_2_42410),
    .O(seg_9_12_sp4_r_v_b_15_38713)
  );
  Span4Mux_h4 t4979 (
    .I(seg_14_9_sp4_v_b_9_53550),
    .O(seg_10_9_sp4_h_r_2_42410)
  );
  CascadeMux t498 (
    .I(net_35552),
    .O(net_35552_cascademuxed)
  );
  LocalMux t4980 (
    .I(seg_9_13_sp4_r_v_b_2_38713),
    .O(seg_9_13_local_g1_2_38983)
  );
  Span4Mux_v4 t4981 (
    .I(seg_10_9_sp4_h_r_2_42410),
    .O(seg_9_13_sp4_r_v_b_2_38713)
  );
  LocalMux t4982 (
    .I(seg_10_13_sp4_v_b_2_38713),
    .O(seg_10_13_local_g1_2_42814)
  );
  Span4Mux_v4 t4983 (
    .I(seg_10_9_sp4_h_r_2_42410),
    .O(seg_10_13_sp4_v_b_2_38713)
  );
  LocalMux t4984 (
    .I(seg_11_17_sp4_h_r_13_43390),
    .O(seg_11_17_local_g0_5_47132)
  );
  Span4Mux_h3 t4985 (
    .I(seg_14_17_sp4_v_b_7_54532),
    .O(seg_11_17_sp4_h_r_13_43390)
  );
  Span4Mux_v4 t4986 (
    .I(seg_14_13_sp4_v_b_11_54044),
    .O(seg_14_17_sp4_v_b_7_54532)
  );
  Span4Mux_v4 t4987 (
    .I(seg_14_9_sp4_v_b_11_53552),
    .O(seg_14_13_sp4_v_b_11_54044)
  );
  LocalMux t4988 (
    .I(seg_9_15_sp4_r_v_b_1_38956),
    .O(seg_9_15_local_g1_1_39228)
  );
  Span4Mux_v4 t4989 (
    .I(seg_10_11_sp4_h_r_1_42653),
    .O(seg_9_15_sp4_r_v_b_1_38956)
  );
  CascadeMux t499 (
    .I(net_35564),
    .O(net_35564_cascademuxed)
  );
  Span4Mux_h4 t4990 (
    .I(seg_14_11_sp4_v_b_1_53788),
    .O(seg_10_11_sp4_h_r_1_42653)
  );
  LocalMux t4991 (
    .I(seg_13_11_sp4_r_v_b_11_53798),
    .O(seg_13_11_local_g2_3_54070)
  );
  LocalMux t4992 (
    .I(seg_14_8_neigh_op_top_0_53764),
    .O(seg_14_8_local_g0_0_57512)
  );
  LocalMux t4993 (
    .I(seg_14_9_lutff_1_out_53765),
    .O(seg_14_9_local_g1_1_57644)
  );
  LocalMux t4994 (
    .I(seg_16_12_sp4_h_r_15_61932),
    .O(seg_16_12_local_g0_7_65672)
  );
  Span4Mux_h1 t4995 (
    .I(seg_15_12_sp4_v_b_8_57750),
    .O(seg_16_12_sp4_h_r_15_61932)
  );
  LocalMux t4996 (
    .I(seg_25_11_sp4_v_b_45_95822),
    .O(seg_25_11_local_g2_5_100171)
  );
  Span4Mux_v1 t4997 (
    .I(seg_25_10_sp4_h_l_45_84047),
    .O(seg_25_11_sp4_v_b_45_95822)
  );
  Sp12to4 t4998 (
    .I(seg_22_10_sp12_h_r_18_54019),
    .O(seg_25_10_sp4_h_l_45_84047)
  );
  LocalMux t4999 (
    .I(seg_25_11_sp4_v_b_41_95818),
    .O(seg_25_11_local_g3_1_100175)
  );
  CascadeMux t50 (
    .I(net_9001),
    .O(net_9001_cascademuxed)
  );
  CascadeMux t500 (
    .I(net_35582),
    .O(net_35582_cascademuxed)
  );
  Span4Mux_v1 t5000 (
    .I(seg_25_10_sp4_h_l_46_84040),
    .O(seg_25_11_sp4_v_b_41_95818)
  );
  Span4Mux_h4 t5001 (
    .I(seg_21_10_sp4_h_l_46_69347),
    .O(seg_25_10_sp4_h_l_46_84040)
  );
  Span4Mux_h4 t5002 (
    .I(seg_17_10_sp4_h_l_38_54027),
    .O(seg_21_10_sp4_h_l_46_69347)
  );
  LocalMux t5003 (
    .I(seg_25_11_sp4_v_b_44_95821),
    .O(seg_25_11_local_g3_4_100178)
  );
  Span4Mux_v1 t5004 (
    .I(seg_25_10_sp4_h_l_41_84043),
    .O(seg_25_11_sp4_v_b_44_95821)
  );
  Span4Mux_h4 t5005 (
    .I(seg_21_10_sp4_h_l_36_69345),
    .O(seg_25_10_sp4_h_l_41_84043)
  );
  Span4Mux_h4 t5006 (
    .I(seg_17_10_sp4_h_l_40_54029),
    .O(seg_21_10_sp4_h_l_36_69345)
  );
  LocalMux t5007 (
    .I(seg_25_12_sp4_v_b_33_95821),
    .O(seg_25_12_local_g2_1_100317)
  );
  Span4Mux_v2 t5008 (
    .I(seg_25_10_sp4_h_l_41_84043),
    .O(seg_25_12_sp4_v_b_33_95821)
  );
  LocalMux t5009 (
    .I(seg_25_11_sp4_v_b_38_95815),
    .O(seg_25_11_local_g3_6_100180)
  );
  Span4Mux_v1 t5010 (
    .I(seg_25_10_sp4_h_l_38_84042),
    .O(seg_25_11_sp4_v_b_38_95815)
  );
  Span4Mux_h4 t5011 (
    .I(seg_21_10_sp4_h_l_38_69349),
    .O(seg_25_10_sp4_h_l_38_84042)
  );
  Span4Mux_h4 t5012 (
    .I(seg_17_10_sp4_h_l_42_54031),
    .O(seg_21_10_sp4_h_l_38_69349)
  );
  LocalMux t5013 (
    .I(seg_25_11_sp4_v_b_39_95816),
    .O(seg_25_11_local_g3_7_100181)
  );
  Span4Mux_v1 t5014 (
    .I(seg_25_10_sp4_h_l_44_84048),
    .O(seg_25_11_sp4_v_b_39_95816)
  );
  Span4Mux_h4 t5015 (
    .I(seg_21_10_sp4_h_l_44_69355),
    .O(seg_25_10_sp4_h_l_44_84048)
  );
  Span4Mux_h4 t5016 (
    .I(seg_17_10_sp4_h_l_44_54033),
    .O(seg_21_10_sp4_h_l_44_69355)
  );
  LocalMux t5017 (
    .I(seg_25_12_sp4_v_b_26_95816),
    .O(seg_25_12_local_g2_2_100318)
  );
  Span4Mux_v2 t5018 (
    .I(seg_25_10_sp4_h_l_44_84048),
    .O(seg_25_12_sp4_v_b_26_95816)
  );
  LocalMux t5019 (
    .I(seg_25_11_sp4_v_b_42_95819),
    .O(seg_25_11_local_g3_2_100176)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t502 (
    .carryinitin(),
    .carryinitout(t501)
  );
  Span4Mux_v1 t5020 (
    .I(seg_25_10_sp4_h_l_42_84046),
    .O(seg_25_11_sp4_v_b_42_95819)
  );
  Span4Mux_h4 t5021 (
    .I(seg_21_10_sp4_h_l_42_69353),
    .O(seg_25_10_sp4_h_l_42_84046)
  );
  Span4Mux_h4 t5022 (
    .I(seg_17_10_sp4_h_l_46_54025),
    .O(seg_21_10_sp4_h_l_42_69353)
  );
  LocalMux t5023 (
    .I(seg_25_12_sp4_v_b_34_95824),
    .O(seg_25_12_local_g3_2_100326)
  );
  Span4Mux_v2 t5024 (
    .I(seg_25_10_sp4_h_l_47_84039),
    .O(seg_25_12_sp4_v_b_34_95824)
  );
  Span4Mux_h4 t5025 (
    .I(seg_21_10_sp4_h_l_42_69353),
    .O(seg_25_10_sp4_h_l_47_84039)
  );
  LocalMux t5026 (
    .I(seg_25_11_sp4_h_r_26_91826),
    .O(seg_25_11_local_g2_2_100168)
  );
  Span4Mux_h2 t5027 (
    .I(seg_23_11_sp4_h_l_43_76905),
    .O(seg_25_11_sp4_h_r_26_91826)
  );
  Span4Mux_h4 t5028 (
    .I(seg_19_11_sp4_h_l_43_61813),
    .O(seg_23_11_sp4_h_l_43_76905)
  );
  Span4Mux_h4 t5029 (
    .I(seg_15_11_sp4_v_b_0_57619),
    .O(seg_19_11_sp4_h_l_43_61813)
  );
  CascadeMux t503 (
    .I(net_37498),
    .O(net_37498_cascademuxed)
  );
  LocalMux t5030 (
    .I(seg_25_12_sp4_h_r_30_91953),
    .O(seg_25_12_local_g3_6_100330)
  );
  Span4Mux_h2 t5031 (
    .I(seg_23_12_sp4_h_l_43_77007),
    .O(seg_25_12_sp4_h_r_30_91953)
  );
  Span4Mux_h4 t5032 (
    .I(seg_19_12_sp4_h_l_38_61933),
    .O(seg_23_12_sp4_h_l_43_77007)
  );
  Span4Mux_h4 t5033 (
    .I(seg_15_12_sp4_v_b_3_57743),
    .O(seg_19_12_sp4_h_l_38_61933)
  );
  LocalMux t5034 (
    .I(seg_25_12_sp4_h_r_25_91946),
    .O(seg_25_12_local_g3_1_100325)
  );
  Span4Mux_h2 t5035 (
    .I(seg_23_12_sp4_h_l_40_77006),
    .O(seg_25_12_sp4_h_r_25_91946)
  );
  Span4Mux_h4 t5036 (
    .I(seg_19_12_sp4_h_l_40_61935),
    .O(seg_23_12_sp4_h_l_40_77006)
  );
  Span4Mux_h4 t5037 (
    .I(seg_15_12_sp4_v_b_5_57745),
    .O(seg_19_12_sp4_h_l_40_61935)
  );
  LocalMux t5038 (
    .I(seg_25_12_sp4_h_r_31_91954),
    .O(seg_25_12_local_g3_7_100331)
  );
  Span4Mux_h2 t5039 (
    .I(seg_23_12_sp4_h_l_42_77008),
    .O(seg_25_12_sp4_h_r_31_91954)
  );
  CascadeMux t504 (
    .I(net_37510),
    .O(net_37510_cascademuxed)
  );
  Span4Mux_h4 t5040 (
    .I(seg_19_12_sp4_h_l_42_61937),
    .O(seg_23_12_sp4_h_l_42_77008)
  );
  Span4Mux_h4 t5041 (
    .I(seg_15_12_sp4_v_b_7_57747),
    .O(seg_19_12_sp4_h_l_42_61937)
  );
  LocalMux t5042 (
    .I(seg_25_12_sp4_h_r_35_91948),
    .O(seg_25_12_local_g2_3_100319)
  );
  Span4Mux_h2 t5043 (
    .I(seg_23_12_sp4_h_l_46_77002),
    .O(seg_25_12_sp4_h_r_35_91948)
  );
  Span4Mux_h4 t5044 (
    .I(seg_19_12_sp4_h_l_46_61931),
    .O(seg_23_12_sp4_h_l_46_77002)
  );
  Span4Mux_h4 t5045 (
    .I(seg_15_12_sp4_v_b_11_57751),
    .O(seg_19_12_sp4_h_l_46_61931)
  );
  LocalMux t5046 (
    .I(seg_14_8_sp4_v_b_32_53674),
    .O(seg_14_8_local_g2_0_57528)
  );
  LocalMux t5047 (
    .I(seg_16_12_sp4_v_b_37_61941),
    .O(seg_16_12_local_g2_5_65686)
  );
  Span4Mux_v1 t5048 (
    .I(seg_16_11_sp4_h_l_37_50314),
    .O(seg_16_12_sp4_v_b_37_61941)
  );
  LocalMux t5049 (
    .I(seg_16_12_sp4_h_r_21_61938),
    .O(seg_16_12_local_g0_5_65670)
  );
  CascadeMux t505 (
    .I(net_37516),
    .O(net_37516_cascademuxed)
  );
  Span4Mux_h1 t5050 (
    .I(seg_15_12_sp4_v_b_2_57744),
    .O(seg_16_12_sp4_h_r_21_61938)
  );
  LocalMux t5051 (
    .I(seg_16_12_sp4_h_r_17_61934),
    .O(seg_16_12_local_g1_1_65674)
  );
  Span4Mux_h1 t5052 (
    .I(seg_15_12_sp4_v_b_4_57746),
    .O(seg_16_12_sp4_h_r_17_61934)
  );
  LocalMux t5053 (
    .I(seg_16_12_sp4_h_r_23_61930),
    .O(seg_16_12_local_g1_7_65680)
  );
  Span4Mux_h1 t5054 (
    .I(seg_15_12_sp4_v_b_10_57752),
    .O(seg_16_12_sp4_h_r_23_61930)
  );
  LocalMux t5055 (
    .I(seg_14_13_neigh_op_bot_4_54137),
    .O(seg_14_13_local_g1_4_58139)
  );
  LocalMux t5056 (
    .I(seg_14_14_sp4_v_b_16_54284),
    .O(seg_14_14_local_g0_0_58250)
  );
  LocalMux t5057 (
    .I(seg_14_10_sp4_v_b_32_53920),
    .O(seg_14_10_local_g2_0_57774)
  );
  LocalMux t5058 (
    .I(seg_15_14_neigh_op_bnl_0_54256),
    .O(seg_15_14_local_g2_0_62096)
  );
  LocalMux t5059 (
    .I(seg_14_13_lutff_1_out_54257),
    .O(seg_14_13_local_g3_1_58152)
  );
  CascadeMux t506 (
    .I(net_37691),
    .O(net_37691_cascademuxed)
  );
  LocalMux t5060 (
    .I(seg_14_13_lutff_3_out_54259),
    .O(seg_14_13_local_g3_3_58154)
  );
  LocalMux t5061 (
    .I(seg_14_14_neigh_op_bot_3_54259),
    .O(seg_14_14_local_g0_3_58253)
  );
  LocalMux t5062 (
    .I(seg_14_13_lutff_4_out_54260),
    .O(seg_14_13_local_g0_4_58131)
  );
  LocalMux t5063 (
    .I(seg_14_13_lutff_6_out_54262),
    .O(seg_14_13_local_g0_6_58133)
  );
  LocalMux t5064 (
    .I(seg_14_14_neigh_op_bot_6_54262),
    .O(seg_14_14_local_g1_6_58264)
  );
  LocalMux t5065 (
    .I(seg_9_13_sp12_h_r_3_35232),
    .O(seg_9_13_local_g1_3_38984)
  );
  LocalMux t5066 (
    .I(seg_14_19_sp12_v_b_0_57482),
    .O(seg_14_19_local_g3_0_58889)
  );
  LocalMux t5067 (
    .I(seg_16_13_sp4_h_r_24_58221),
    .O(seg_16_13_local_g3_0_65812)
  );
  LocalMux t5068 (
    .I(seg_16_13_sp4_h_r_34_58223),
    .O(seg_16_13_local_g2_2_65806)
  );
  LocalMux t5069 (
    .I(seg_9_14_sp4_v_b_46_35381),
    .O(seg_9_14_local_g2_6_39118)
  );
  CascadeMux t507 (
    .I(net_37814),
    .O(net_37814_cascademuxed)
  );
  Span4Mux_v1 t5070 (
    .I(seg_9_13_sp4_h_r_11_39070),
    .O(seg_9_14_sp4_v_b_46_35381)
  );
  Span4Mux_h4 t5071 (
    .I(seg_13_13_sp4_h_r_3_54396),
    .O(seg_9_13_sp4_h_r_11_39070)
  );
  LocalMux t5072 (
    .I(seg_10_14_sp4_r_v_b_42_43039),
    .O(seg_10_14_local_g3_2_42953)
  );
  Span4Mux_v1 t5073 (
    .I(seg_11_13_sp4_h_r_1_46730),
    .O(seg_10_14_sp4_r_v_b_42_43039)
  );
  LocalMux t5074 (
    .I(seg_11_13_sp4_h_r_1_46730),
    .O(seg_11_13_local_g1_1_46644)
  );
  LocalMux t5075 (
    .I(seg_10_14_sp4_r_v_b_40_43037),
    .O(seg_10_14_local_g3_0_42951)
  );
  Span4Mux_v1 t5076 (
    .I(seg_11_13_sp4_h_r_11_46732),
    .O(seg_10_14_sp4_r_v_b_40_43037)
  );
  LocalMux t5077 (
    .I(seg_10_15_sp4_r_v_b_29_43037),
    .O(seg_10_15_local_g1_5_43063)
  );
  Span4Mux_v2 t5078 (
    .I(seg_11_13_sp4_h_r_11_46732),
    .O(seg_10_15_sp4_r_v_b_29_43037)
  );
  LocalMux t5079 (
    .I(seg_11_14_sp4_h_r_8_46862),
    .O(seg_11_14_local_g0_0_46758)
  );
  CascadeMux t508 (
    .I(net_37901),
    .O(net_37901_cascademuxed)
  );
  Span4Mux_h4 t5080 (
    .I(seg_15_14_sp4_v_b_8_57996),
    .O(seg_11_14_sp4_h_r_8_46862)
  );
  LocalMux t5081 (
    .I(seg_14_15_sp4_r_v_b_5_58114),
    .O(seg_14_15_local_g1_5_58386)
  );
  LocalMux t5082 (
    .I(seg_9_15_sp4_h_r_27_31656),
    .O(seg_9_15_local_g3_3_39246)
  );
  Span4Mux_h2 t5083 (
    .I(seg_11_15_sp4_h_r_0_46975),
    .O(seg_9_15_sp4_h_r_27_31656)
  );
  Span4Mux_h4 t5084 (
    .I(seg_15_15_sp4_v_b_7_58116),
    .O(seg_11_15_sp4_h_r_0_46975)
  );
  LocalMux t5085 (
    .I(seg_14_15_sp4_r_v_b_15_58236),
    .O(seg_14_15_local_g2_7_58396)
  );
  LocalMux t5086 (
    .I(seg_14_19_sp4_r_v_b_23_58736),
    .O(seg_14_19_local_g3_7_58896)
  );
  Span4Mux_v3 t5087 (
    .I(seg_15_16_sp4_v_b_2_58236),
    .O(seg_14_19_sp4_r_v_b_23_58736)
  );
  LocalMux t5088 (
    .I(seg_14_14_lutff_0_out_54379),
    .O(seg_14_14_local_g3_0_58274)
  );
  LocalMux t5089 (
    .I(seg_14_15_neigh_op_bot_0_54379),
    .O(seg_14_15_local_g0_0_58373)
  );
  CascadeMux t509 (
    .I(net_37937),
    .O(net_37937_cascademuxed)
  );
  LocalMux t5090 (
    .I(seg_14_14_lutff_2_out_54381),
    .O(seg_14_14_local_g2_2_58268)
  );
  LocalMux t5091 (
    .I(seg_14_15_neigh_op_bot_2_54381),
    .O(seg_14_15_local_g0_2_58375)
  );
  LocalMux t5092 (
    .I(seg_14_14_lutff_4_out_54383),
    .O(seg_14_14_local_g2_4_58270)
  );
  LocalMux t5093 (
    .I(seg_14_15_neigh_op_bot_4_54383),
    .O(seg_14_15_local_g1_4_58385)
  );
  LocalMux t5094 (
    .I(seg_14_15_neigh_op_bot_5_54384),
    .O(seg_14_15_local_g0_5_58378)
  );
  LocalMux t5095 (
    .I(seg_14_15_neigh_op_bot_6_54385),
    .O(seg_14_15_local_g1_6_58387)
  );
  LocalMux t5096 (
    .I(seg_14_14_lutff_7_out_54386),
    .O(seg_14_14_local_g2_7_58273)
  );
  LocalMux t5097 (
    .I(seg_14_15_neigh_op_bot_7_54386),
    .O(seg_14_15_local_g1_7_58388)
  );
  LocalMux t5098 (
    .I(seg_14_19_sp12_v_b_3_57605),
    .O(seg_14_19_local_g3_3_58892)
  );
  LocalMux t5099 (
    .I(seg_18_12_sp4_v_b_34_69490),
    .O(seg_18_12_local_g3_2_73353)
  );
  CascadeMux t51 (
    .I(net_9154),
    .O(net_9154_cascademuxed)
  );
  CascadeMux t510 (
    .I(net_38024),
    .O(net_38024_cascademuxed)
  );
  Span4Mux_v2 t5100 (
    .I(seg_18_14_sp4_h_l_47_58346),
    .O(seg_18_12_sp4_v_b_34_69490)
  );
  LocalMux t5101 (
    .I(seg_18_14_sp4_h_r_26_66009),
    .O(seg_18_14_local_g3_2_73599)
  );
  Span4Mux_h2 t5102 (
    .I(seg_16_14_sp4_h_l_43_50691),
    .O(seg_18_14_sp4_h_r_26_66009)
  );
  LocalMux t5103 (
    .I(seg_18_13_sp4_v_b_17_69484),
    .O(seg_18_13_local_g0_1_73451)
  );
  Span4Mux_v1 t5104 (
    .I(seg_18_14_sp4_h_l_41_58350),
    .O(seg_18_13_sp4_v_b_17_69484)
  );
  LocalMux t5105 (
    .I(seg_18_14_sp4_h_r_11_73670),
    .O(seg_18_14_local_g1_3_73584)
  );
  Span4Mux_h0 t5106 (
    .I(seg_18_14_sp4_h_l_45_58354),
    .O(seg_18_14_sp4_h_r_11_73670)
  );
  LocalMux t5107 (
    .I(seg_15_12_sp4_v_b_25_57987),
    .O(seg_15_12_local_g2_1_61851)
  );
  LocalMux t5108 (
    .I(seg_15_16_sp4_v_b_9_58241),
    .O(seg_15_16_local_g0_1_62327)
  );
  LocalMux t5109 (
    .I(seg_15_16_sp4_v_b_13_58357),
    .O(seg_15_16_local_g0_5_62331)
  );
  CascadeMux t511 (
    .I(net_38060),
    .O(net_38060_cascademuxed)
  );
  LocalMux t5110 (
    .I(seg_15_16_sp4_v_b_17_58361),
    .O(seg_15_16_local_g1_1_62335)
  );
  LocalMux t5111 (
    .I(seg_15_16_sp4_v_b_19_58363),
    .O(seg_15_16_local_g1_3_62337)
  );
  LocalMux t5112 (
    .I(seg_16_17_sp4_h_r_19_62551),
    .O(seg_16_17_local_g0_3_66283)
  );
  Span4Mux_h1 t5113 (
    .I(seg_15_17_sp4_v_b_6_58363),
    .O(seg_16_17_sp4_h_r_19_62551)
  );
  LocalMux t5114 (
    .I(seg_15_16_sp4_v_b_23_58367),
    .O(seg_15_16_local_g0_7_62333)
  );
  LocalMux t5115 (
    .I(seg_14_16_neigh_op_bot_0_54502),
    .O(seg_14_16_local_g1_0_58504)
  );
  LocalMux t5116 (
    .I(seg_13_14_neigh_op_tnr_2_54504),
    .O(seg_13_14_local_g2_2_54438)
  );
  LocalMux t5117 (
    .I(seg_13_15_neigh_op_rgt_2_54504),
    .O(seg_13_15_local_g2_2_54561)
  );
  LocalMux t5118 (
    .I(seg_14_16_neigh_op_bot_3_54505),
    .O(seg_14_16_local_g0_3_58499)
  );
  LocalMux t5119 (
    .I(seg_14_15_lutff_4_out_54506),
    .O(seg_14_15_local_g2_4_58393)
  );
  CascadeMux t512 (
    .I(net_38276),
    .O(net_38276_cascademuxed)
  );
  LocalMux t5120 (
    .I(seg_14_16_neigh_op_bot_5_54507),
    .O(seg_14_16_local_g0_5_58501)
  );
  LocalMux t5121 (
    .I(seg_14_16_neigh_op_bot_6_54508),
    .O(seg_14_16_local_g1_6_58510)
  );
  LocalMux t5122 (
    .I(seg_14_16_neigh_op_bot_7_54509),
    .O(seg_14_16_local_g1_7_58511)
  );
  LocalMux t5123 (
    .I(seg_14_19_sp12_v_b_10_58096),
    .O(seg_14_19_local_g2_2_58883)
  );
  LocalMux t5124 (
    .I(seg_12_15_sp4_h_r_12_46976),
    .O(seg_12_15_local_g1_4_50724)
  );
  LocalMux t5125 (
    .I(seg_14_13_sp4_v_b_32_54289),
    .O(seg_14_13_local_g3_0_58151)
  );
  LocalMux t5126 (
    .I(seg_16_16_sp4_h_r_38_54765),
    .O(seg_16_16_local_g3_6_66187)
  );
  LocalMux t5127 (
    .I(seg_16_16_sp4_h_r_3_66256),
    .O(seg_16_16_local_g0_3_66160)
  );
  Span4Mux_h0 t5128 (
    .I(seg_16_16_sp4_h_l_37_50929),
    .O(seg_16_16_sp4_h_r_3_66256)
  );
  LocalMux t5129 (
    .I(seg_16_16_sp4_h_r_28_58596),
    .O(seg_16_16_local_g3_4_66185)
  );
  CascadeMux t513 (
    .I(net_38294),
    .O(net_38294_cascademuxed)
  );
  LocalMux t5130 (
    .I(seg_16_16_sp4_h_r_22_62423),
    .O(seg_16_16_local_g1_6_66171)
  );
  Span4Mux_h1 t5131 (
    .I(seg_15_16_sp4_v_b_11_58243),
    .O(seg_16_16_sp4_h_r_22_62423)
  );
  LocalMux t5132 (
    .I(seg_14_18_sp4_r_v_b_15_58605),
    .O(seg_14_18_local_g2_7_58765)
  );
  LocalMux t5133 (
    .I(seg_14_18_sp4_v_b_20_54780),
    .O(seg_14_18_local_g1_4_58754)
  );
  LocalMux t5134 (
    .I(seg_14_17_lutff_2_out_54750),
    .O(seg_14_17_local_g0_2_58621)
  );
  LocalMux t5135 (
    .I(seg_14_17_lutff_3_out_54751),
    .O(seg_14_17_local_g3_3_58646)
  );
  LocalMux t5136 (
    .I(seg_14_18_neigh_op_bot_5_54753),
    .O(seg_14_18_local_g0_5_58747)
  );
  LocalMux t5137 (
    .I(seg_14_18_neigh_op_bot_6_54754),
    .O(seg_14_18_local_g1_6_58756)
  );
  LocalMux t5138 (
    .I(seg_14_16_neigh_op_top_7_54755),
    .O(seg_14_16_local_g0_7_58503)
  );
  LocalMux t5139 (
    .I(seg_16_17_sp4_h_r_24_58713),
    .O(seg_16_17_local_g3_0_66304)
  );
  CascadeMux t514 (
    .I(net_38312),
    .O(net_38312_cascademuxed)
  );
  LocalMux t5140 (
    .I(seg_17_17_sp4_h_r_39_58717),
    .O(seg_17_17_local_g2_7_70134)
  );
  LocalMux t5141 (
    .I(seg_17_14_sp4_h_r_30_62182),
    .O(seg_17_14_local_g2_6_69764)
  );
  Span4Mux_h2 t5142 (
    .I(seg_15_14_sp4_v_t_43_58486),
    .O(seg_17_14_sp4_h_r_30_62182)
  );
  LocalMux t5143 (
    .I(seg_17_13_sp4_h_r_27_62056),
    .O(seg_17_13_local_g2_3_69638)
  );
  Span4Mux_h2 t5144 (
    .I(seg_15_13_sp4_v_t_38_58358),
    .O(seg_17_13_sp4_h_r_27_62056)
  );
  LocalMux t5145 (
    .I(seg_14_18_lutff_0_out_54871),
    .O(seg_14_18_local_g1_0_58750)
  );
  LocalMux t5146 (
    .I(seg_14_17_neigh_op_top_1_54872),
    .O(seg_14_17_local_g0_1_58620)
  );
  LocalMux t5147 (
    .I(seg_15_17_neigh_op_tnl_1_54872),
    .O(seg_15_17_local_g2_1_62466)
  );
  LocalMux t5148 (
    .I(seg_14_18_lutff_3_out_54874),
    .O(seg_14_18_local_g3_3_58769)
  );
  LocalMux t5149 (
    .I(seg_15_17_neigh_op_tnl_5_54876),
    .O(seg_15_17_local_g2_5_62470)
  );
  CascadeMux t515 (
    .I(net_38393),
    .O(net_38393_cascademuxed)
  );
  LocalMux t5150 (
    .I(seg_14_17_neigh_op_top_7_54878),
    .O(seg_14_17_local_g0_7_58626)
  );
  LocalMux t5151 (
    .I(seg_15_17_neigh_op_tnl_7_54878),
    .O(seg_15_17_local_g3_7_62480)
  );
  LocalMux t5152 (
    .I(seg_15_16_sp4_v_b_35_58489),
    .O(seg_15_16_local_g2_3_62345)
  );
  LocalMux t5153 (
    .I(seg_15_16_sp4_v_b_37_58603),
    .O(seg_15_16_local_g3_5_62355)
  );
  LocalMux t5154 (
    .I(seg_14_16_sp4_r_v_b_27_58481),
    .O(seg_14_16_local_g1_3_58507)
  );
  LocalMux t5155 (
    .I(seg_15_16_sp4_v_b_27_58481),
    .O(seg_15_16_local_g3_3_62353)
  );
  LocalMux t5156 (
    .I(seg_14_16_sp4_r_v_b_29_58483),
    .O(seg_14_16_local_g1_5_58509)
  );
  LocalMux t5157 (
    .I(seg_15_16_sp4_v_b_29_58483),
    .O(seg_15_16_local_g2_5_62347)
  );
  LocalMux t5158 (
    .I(seg_14_16_sp4_v_b_34_54660),
    .O(seg_14_16_local_g2_2_58514)
  );
  LocalMux t5159 (
    .I(seg_14_16_sp4_v_b_36_54772),
    .O(seg_14_16_local_g2_4_58516)
  );
  CascadeMux t516 (
    .I(net_38399),
    .O(net_38399_cascademuxed)
  );
  LocalMux t5160 (
    .I(seg_14_19_lutff_3_out_54997),
    .O(seg_14_19_local_g2_3_58884)
  );
  LocalMux t5161 (
    .I(seg_12_16_sp4_h_r_29_43274),
    .O(seg_12_16_local_g2_5_50856)
  );
  Span4Mux_h2 t5162 (
    .I(seg_14_16_sp4_v_t_46_54905),
    .O(seg_12_16_sp4_h_r_29_43274)
  );
  LocalMux t5163 (
    .I(seg_13_16_sp4_h_r_40_43274),
    .O(seg_13_16_local_g2_0_54682)
  );
  Span4Mux_h1 t5164 (
    .I(seg_14_16_sp4_v_t_46_54905),
    .O(seg_13_16_sp4_h_r_40_43274)
  );
  LocalMux t5165 (
    .I(seg_14_15_sp4_v_b_15_54406),
    .O(seg_14_15_local_g0_7_58380)
  );
  Span4Mux_v1 t5166 (
    .I(seg_14_16_sp4_v_t_46_54905),
    .O(seg_14_15_sp4_v_b_15_54406)
  );
  LocalMux t5167 (
    .I(seg_3_2_sp4_v_b_22_11410),
    .O(seg_3_2_local_g1_6_15279)
  );
  Span4Mux_v1 t5168 (
    .I(seg_3_3_sp4_h_r_11_15485),
    .O(seg_3_2_sp4_v_b_22_11410)
  );
  Span4Mux_h4 t5169 (
    .I(seg_7_3_sp4_h_r_3_30180),
    .O(seg_3_3_sp4_h_r_11_15485)
  );
  CascadeMux t517 (
    .I(net_38411),
    .O(net_38411_cascademuxed)
  );
  Span4Mux_h4 t5170 (
    .I(seg_11_3_sp4_h_r_0_45499),
    .O(seg_7_3_sp4_h_r_3_30180)
  );
  Span4Mux_h4 t5171 (
    .I(seg_15_3_sp4_v_b_0_56738),
    .O(seg_11_3_sp4_h_r_0_45499)
  );
  LocalMux t5172 (
    .I(seg_3_3_sp4_h_r_11_15485),
    .O(seg_3_3_local_g0_3_15391)
  );
  LocalMux t5173 (
    .I(seg_4_3_sp4_h_r_22_15485),
    .O(seg_4_3_local_g1_6_19233)
  );
  Span4Mux_h3 t5174 (
    .I(seg_7_3_sp4_h_r_3_30180),
    .O(seg_4_3_sp4_h_r_22_15485)
  );
  LocalMux t5175 (
    .I(seg_15_6_sp4_v_b_31_57255),
    .O(seg_15_6_local_g3_7_61127)
  );
  Span4Mux_v2 t5176 (
    .I(seg_15_4_sp4_v_b_4_56757),
    .O(seg_15_6_sp4_v_b_31_57255)
  );
  LocalMux t5177 (
    .I(seg_16_4_neigh_op_bnl_2_56858),
    .O(seg_16_4_local_g2_2_64699)
  );
  LocalMux t5178 (
    .I(seg_13_3_sp4_h_r_16_49337),
    .O(seg_13_3_local_g0_0_53067)
  );
  LocalMux t5179 (
    .I(seg_15_4_lutff_0_out_56979),
    .O(seg_15_4_local_g0_0_60850)
  );
  CascadeMux t518 (
    .I(net_38423),
    .O(net_38423_cascademuxed)
  );
  LocalMux t5180 (
    .I(seg_15_3_neigh_op_top_2_56981),
    .O(seg_15_3_local_g0_2_60729)
  );
  LocalMux t5181 (
    .I(seg_16_4_neigh_op_lft_7_56986),
    .O(seg_16_4_local_g0_7_64688)
  );
  LocalMux t5182 (
    .I(seg_25_6_sp4_v_b_32_94988),
    .O(seg_25_6_local_g3_0_99394)
  );
  Span4Mux_v2 t5183 (
    .I(seg_25_4_sp4_h_l_45_83309),
    .O(seg_25_6_sp4_v_b_32_94988)
  );
  Span4Mux_h4 t5184 (
    .I(seg_21_4_sp4_h_l_37_68606),
    .O(seg_25_4_sp4_h_l_45_83309)
  );
  Span4Mux_h4 t5185 (
    .I(seg_17_4_sp4_h_l_37_53284),
    .O(seg_21_4_sp4_h_l_37_68606)
  );
  LocalMux t5186 (
    .I(seg_25_6_sp4_v_b_34_94990),
    .O(seg_25_6_local_g3_2_99396)
  );
  Span4Mux_v2 t5187 (
    .I(seg_25_4_sp4_h_l_47_83301),
    .O(seg_25_6_sp4_v_b_34_94990)
  );
  Span4Mux_h4 t5188 (
    .I(seg_21_4_sp4_h_l_39_68610),
    .O(seg_25_4_sp4_h_l_47_83301)
  );
  Span4Mux_h4 t5189 (
    .I(seg_17_4_sp4_h_l_39_53288),
    .O(seg_21_4_sp4_h_l_39_68610)
  );
  CascadeMux t519 (
    .I(net_38429),
    .O(net_38429_cascademuxed)
  );
  LocalMux t5190 (
    .I(seg_25_7_sp4_v_b_18_94985),
    .O(seg_25_7_local_g1_2_99530)
  );
  Span4Mux_v3 t5191 (
    .I(seg_25_4_sp4_h_l_39_83303),
    .O(seg_25_7_sp4_v_b_18_94985)
  );
  Span4Mux_h4 t5192 (
    .I(seg_21_4_sp4_h_l_39_68610),
    .O(seg_25_4_sp4_h_l_39_83303)
  );
  LocalMux t5193 (
    .I(seg_25_6_sp4_v_b_26_94982),
    .O(seg_25_6_local_g2_2_99388)
  );
  Span4Mux_v2 t5194 (
    .I(seg_25_4_sp4_h_l_44_83310),
    .O(seg_25_6_sp4_v_b_26_94982)
  );
  Span4Mux_h4 t5195 (
    .I(seg_21_4_sp4_h_l_43_68614),
    .O(seg_25_4_sp4_h_l_44_83310)
  );
  Span4Mux_h4 t5196 (
    .I(seg_17_4_sp4_h_l_47_53286),
    .O(seg_21_4_sp4_h_l_43_68614)
  );
  LocalMux t5197 (
    .I(seg_25_7_sp4_v_b_15_94982),
    .O(seg_25_7_local_g1_7_99535)
  );
  Span4Mux_v3 t5198 (
    .I(seg_25_4_sp4_h_l_44_83310),
    .O(seg_25_7_sp4_v_b_15_94982)
  );
  LocalMux t5199 (
    .I(seg_25_6_sp4_v_b_27_94981),
    .O(seg_25_6_local_g2_3_99389)
  );
  CascadeMux t52 (
    .I(net_9289),
    .O(net_9289_cascademuxed)
  );
  CascadeMux t520 (
    .I(net_38435),
    .O(net_38435_cascademuxed)
  );
  Span4Mux_v2 t5200 (
    .I(seg_25_4_sp4_v_b_3_90450),
    .O(seg_25_6_sp4_v_b_27_94981)
  );
  IoSpan4Mux t5201 (
    .I(seg_23_0_span4_vert_37_86768),
    .O(seg_25_4_sp4_v_b_3_90450)
  );
  Span4Mux_v4 t5202 (
    .I(seg_23_4_sp4_h_l_43_76191),
    .O(seg_23_0_span4_vert_37_86768)
  );
  Span4Mux_h4 t5203 (
    .I(seg_19_4_sp4_h_l_43_60952),
    .O(seg_23_4_sp4_h_l_43_76191)
  );
  LocalMux t5204 (
    .I(seg_25_6_sp4_h_r_16_95113),
    .O(seg_25_6_local_g0_0_99370)
  );
  Span4Mux_h1 t5205 (
    .I(seg_24_6_sp4_h_l_40_79721),
    .O(seg_25_6_sp4_h_r_16_95113)
  );
  Span4Mux_h4 t5206 (
    .I(seg_20_6_sp4_h_l_40_65028),
    .O(seg_24_6_sp4_h_l_40_79721)
  );
  Span4Mux_h4 t5207 (
    .I(seg_16_6_sp4_v_b_5_60837),
    .O(seg_20_6_sp4_h_l_40_65028)
  );
  LocalMux t5208 (
    .I(seg_25_7_sp4_h_r_17_95251),
    .O(seg_25_7_local_g0_1_99521)
  );
  Span4Mux_h1 t5209 (
    .I(seg_24_7_sp4_h_l_41_79843),
    .O(seg_25_7_sp4_h_r_17_95251)
  );
  CascadeMux t521 (
    .I(net_38522),
    .O(net_38522_cascademuxed)
  );
  Span4Mux_h4 t5210 (
    .I(seg_20_7_sp4_h_l_45_65154),
    .O(seg_24_7_sp4_h_l_41_79843)
  );
  Span4Mux_h4 t5211 (
    .I(seg_16_7_sp4_v_b_2_60959),
    .O(seg_20_7_sp4_h_l_45_65154)
  );
  LocalMux t5212 (
    .I(seg_25_7_sp4_h_r_23_95247),
    .O(seg_25_7_local_g0_7_99527)
  );
  Span4Mux_h1 t5213 (
    .I(seg_24_7_sp4_h_l_47_79839),
    .O(seg_25_7_sp4_h_r_23_95247)
  );
  Span4Mux_h4 t5214 (
    .I(seg_20_7_sp4_h_l_47_65146),
    .O(seg_24_7_sp4_h_l_47_79839)
  );
  Span4Mux_h4 t5215 (
    .I(seg_16_7_sp4_v_b_4_60961),
    .O(seg_20_7_sp4_h_l_47_65146)
  );
  LocalMux t5216 (
    .I(seg_25_7_sp4_h_r_33_91341),
    .O(seg_25_7_local_g3_1_99545)
  );
  Span4Mux_h2 t5217 (
    .I(seg_23_7_sp4_h_l_43_76497),
    .O(seg_25_7_sp4_h_r_33_91341)
  );
  Span4Mux_h4 t5218 (
    .I(seg_19_7_sp4_h_l_38_61318),
    .O(seg_23_7_sp4_h_l_43_76497)
  );
  Span4Mux_h4 t5219 (
    .I(seg_15_7_sp4_v_b_9_57134),
    .O(seg_19_7_sp4_h_l_38_61318)
  );
  CascadeMux t522 (
    .I(net_38528),
    .O(net_38528_cascademuxed)
  );
  LocalMux t5220 (
    .I(seg_25_7_sp12_h_r_20_61309),
    .O(seg_25_7_local_g1_4_99532)
  );
  Span12Mux_h10 t5221 (
    .I(seg_15_7_sp12_v_b_0_60411),
    .O(seg_25_7_sp12_h_r_20_61309)
  );
  LocalMux t5222 (
    .I(seg_25_6_sp4_v_b_45_95127),
    .O(seg_25_6_local_g2_5_99391)
  );
  Span4Mux_v1 t5223 (
    .I(seg_25_5_sp4_h_l_45_83432),
    .O(seg_25_6_sp4_v_b_45_95127)
  );
  Span4Mux_h4 t5224 (
    .I(seg_21_5_sp4_h_l_37_68729),
    .O(seg_25_5_sp4_h_l_45_83432)
  );
  Span4Mux_h4 t5225 (
    .I(seg_17_5_sp4_h_l_37_53407),
    .O(seg_21_5_sp4_h_l_37_68729)
  );
  LocalMux t5226 (
    .I(seg_25_7_sp4_v_b_32_95127),
    .O(seg_25_7_local_g3_0_99544)
  );
  Span4Mux_v2 t5227 (
    .I(seg_25_5_sp4_h_l_45_83432),
    .O(seg_25_7_sp4_v_b_32_95127)
  );
  LocalMux t5228 (
    .I(seg_25_6_sp4_v_b_47_95129),
    .O(seg_25_6_local_g3_7_99401)
  );
  Span4Mux_v1 t5229 (
    .I(seg_25_5_sp4_h_l_40_83429),
    .O(seg_25_6_sp4_v_b_47_95129)
  );
  CascadeMux t523 (
    .I(net_38639),
    .O(net_38639_cascademuxed)
  );
  Span4Mux_h4 t5230 (
    .I(seg_21_5_sp4_h_l_39_68733),
    .O(seg_25_5_sp4_h_l_40_83429)
  );
  Span4Mux_h4 t5231 (
    .I(seg_17_5_sp4_h_l_39_53411),
    .O(seg_21_5_sp4_h_l_39_68733)
  );
  LocalMux t5232 (
    .I(seg_25_7_sp4_v_b_29_95122),
    .O(seg_25_7_local_g3_5_99549)
  );
  Span4Mux_v2 t5233 (
    .I(seg_25_5_sp4_h_l_40_83429),
    .O(seg_25_7_sp4_v_b_29_95122)
  );
  LocalMux t5234 (
    .I(seg_25_6_sp4_v_b_37_95119),
    .O(seg_25_6_local_g3_5_99399)
  );
  Span4Mux_v1 t5235 (
    .I(seg_25_5_sp4_h_l_37_83422),
    .O(seg_25_6_sp4_v_b_37_95119)
  );
  Span4Mux_h4 t5236 (
    .I(seg_21_5_sp4_h_l_44_68740),
    .O(seg_25_5_sp4_h_l_37_83422)
  );
  Span4Mux_h4 t5237 (
    .I(seg_17_5_sp4_h_l_43_53415),
    .O(seg_21_5_sp4_h_l_44_68740)
  );
  LocalMux t5238 (
    .I(seg_25_7_sp4_v_b_24_95119),
    .O(seg_25_7_local_g2_0_99536)
  );
  Span4Mux_v2 t5239 (
    .I(seg_25_5_sp4_h_l_37_83422),
    .O(seg_25_7_sp4_v_b_24_95119)
  );
  CascadeMux t524 (
    .I(net_38675),
    .O(net_38675_cascademuxed)
  );
  LocalMux t5240 (
    .I(seg_25_6_sp4_h_r_13_95106),
    .O(seg_25_6_local_g1_5_99383)
  );
  Span4Mux_h1 t5241 (
    .I(seg_24_6_sp4_h_l_44_79725),
    .O(seg_25_6_sp4_h_r_13_95106)
  );
  Span4Mux_h4 t5242 (
    .I(seg_20_6_sp4_h_l_43_65029),
    .O(seg_24_6_sp4_h_l_44_79725)
  );
  Span4Mux_h4 t5243 (
    .I(seg_16_6_sp4_v_b_0_60834),
    .O(seg_20_6_sp4_h_l_43_65029)
  );
  LocalMux t5244 (
    .I(seg_25_6_sp4_h_r_18_95115),
    .O(seg_25_6_local_g1_2_99380)
  );
  Span4Mux_h1 t5245 (
    .I(seg_24_6_sp4_h_l_46_79717),
    .O(seg_25_6_sp4_h_r_18_95115)
  );
  Span4Mux_h4 t5246 (
    .I(seg_20_6_sp4_h_l_45_65031),
    .O(seg_24_6_sp4_h_l_46_79717)
  );
  Span4Mux_h4 t5247 (
    .I(seg_16_6_sp4_v_b_8_60842),
    .O(seg_20_6_sp4_h_l_45_65031)
  );
  LocalMux t5248 (
    .I(seg_25_6_sp4_h_r_23_95108),
    .O(seg_25_6_local_g1_7_99385)
  );
  Span4Mux_h1 t5249 (
    .I(seg_24_6_sp4_h_l_42_79723),
    .O(seg_25_6_sp4_h_r_23_95108)
  );
  CascadeMux t525 (
    .I(net_38891),
    .O(net_38891_cascademuxed)
  );
  Span4Mux_h4 t5250 (
    .I(seg_20_6_sp4_h_l_41_65027),
    .O(seg_24_6_sp4_h_l_42_79723)
  );
  Span4Mux_h4 t5251 (
    .I(seg_16_6_sp4_v_b_10_60844),
    .O(seg_20_6_sp4_h_l_41_65027)
  );
  LocalMux t5252 (
    .I(seg_25_7_sp4_v_b_1_94840),
    .O(seg_25_7_local_g1_1_99529)
  );
  Span4Mux_v4 t5253 (
    .I(seg_25_3_sp4_v_b_10_94273),
    .O(seg_25_7_sp4_v_b_1_94840)
  );
  IoSpan4Mux t5254 (
    .I(seg_24_0_span4_vert_13_90573),
    .O(seg_25_3_sp4_v_b_10_94273)
  );
  Span4Mux_v2 t5255 (
    .I(seg_24_2_sp4_h_l_43_79230),
    .O(seg_24_0_span4_vert_13_90573)
  );
  Span4Mux_h4 t5256 (
    .I(seg_20_2_sp4_h_l_47_64531),
    .O(seg_24_2_sp4_h_l_43_79230)
  );
  Span4Mux_h4 t5257 (
    .I(seg_16_2_sp4_v_t_47_60844),
    .O(seg_20_2_sp4_h_l_47_64531)
  );
  LocalMux t5258 (
    .I(seg_25_7_sp4_h_r_21_95255),
    .O(seg_25_7_local_g1_5_99533)
  );
  Span4Mux_h1 t5259 (
    .I(seg_24_7_sp4_h_l_40_79844),
    .O(seg_25_7_sp4_h_r_21_95255)
  );
  CascadeMux t526 (
    .I(net_39026),
    .O(net_39026_cascademuxed)
  );
  Span4Mux_h4 t5260 (
    .I(seg_20_7_sp4_h_l_40_65151),
    .O(seg_24_7_sp4_h_l_40_79844)
  );
  Span4Mux_h4 t5261 (
    .I(seg_16_7_sp4_v_b_5_60960),
    .O(seg_20_7_sp4_h_l_40_65151)
  );
  LocalMux t5262 (
    .I(seg_25_7_sp4_h_r_19_95253),
    .O(seg_25_7_local_g0_3_99523)
  );
  Span4Mux_h1 t5263 (
    .I(seg_24_7_sp4_h_l_38_79842),
    .O(seg_25_7_sp4_h_r_19_95253)
  );
  Span4Mux_h4 t5264 (
    .I(seg_20_7_sp4_h_l_38_65149),
    .O(seg_24_7_sp4_h_l_38_79842)
  );
  Span4Mux_h4 t5265 (
    .I(seg_16_7_sp4_v_b_9_60964),
    .O(seg_20_7_sp4_h_l_38_65149)
  );
  LocalMux t5266 (
    .I(seg_25_6_sp4_h_r_28_91213),
    .O(seg_25_6_local_g3_4_99398)
  );
  Span4Mux_h2 t5267 (
    .I(seg_23_6_sp4_h_l_36_76388),
    .O(seg_25_6_sp4_h_r_28_91213)
  );
  Span4Mux_h4 t5268 (
    .I(seg_19_6_sp4_h_l_40_61197),
    .O(seg_23_6_sp4_h_l_36_76388)
  );
  Span4Mux_h4 t5269 (
    .I(seg_15_6_sp4_v_b_5_57007),
    .O(seg_19_6_sp4_h_l_40_61197)
  );
  CascadeMux t527 (
    .I(net_39044),
    .O(net_39044_cascademuxed)
  );
  LocalMux t5270 (
    .I(seg_25_6_sp4_h_r_25_91208),
    .O(seg_25_6_local_g3_1_99395)
  );
  Span4Mux_h2 t5271 (
    .I(seg_23_6_sp4_h_l_47_76389),
    .O(seg_25_6_sp4_h_r_25_91208)
  );
  Span4Mux_h4 t5272 (
    .I(seg_19_6_sp4_h_l_42_61199),
    .O(seg_23_6_sp4_h_l_47_76389)
  );
  Span4Mux_h4 t5273 (
    .I(seg_15_6_sp4_v_b_7_57009),
    .O(seg_19_6_sp4_h_l_42_61199)
  );
  LocalMux t5274 (
    .I(seg_25_7_sp4_h_r_27_91335),
    .O(seg_25_7_local_g3_3_99547)
  );
  Span4Mux_h2 t5275 (
    .I(seg_23_7_sp4_h_l_42_76498),
    .O(seg_25_7_sp4_h_r_27_91335)
  );
  Span4Mux_h4 t5276 (
    .I(seg_19_7_sp4_h_l_41_61319),
    .O(seg_23_7_sp4_h_l_42_76498)
  );
  Span4Mux_h4 t5277 (
    .I(seg_15_7_sp4_v_b_10_57137),
    .O(seg_19_7_sp4_h_l_41_61319)
  );
  LocalMux t5278 (
    .I(seg_14_6_neigh_op_rgt_0_57225),
    .O(seg_14_6_local_g2_0_57282)
  );
  LocalMux t5279 (
    .I(seg_14_6_neigh_op_rgt_4_57229),
    .O(seg_14_6_local_g3_4_57294)
  );
  CascadeMux t528 (
    .I(net_39131),
    .O(net_39131_cascademuxed)
  );
  LocalMux t5280 (
    .I(seg_15_7_neigh_op_bot_7_57232),
    .O(seg_15_7_local_g1_7_61234)
  );
  LocalMux t5281 (
    .I(seg_11_9_sp4_v_b_23_42183),
    .O(seg_11_9_local_g1_7_46158)
  );
  Span4Mux_v3 t5282 (
    .I(seg_11_6_sp4_h_r_10_45870),
    .O(seg_11_9_sp4_v_b_23_42183)
  );
  Span4Mux_h4 t5283 (
    .I(seg_15_6_sp4_h_r_2_61194),
    .O(seg_11_6_sp4_h_r_10_45870)
  );
  LocalMux t5284 (
    .I(seg_12_4_sp4_v_b_32_45520),
    .O(seg_12_4_local_g2_0_49375)
  );
  Span4Mux_v2 t5285 (
    .I(seg_12_6_sp4_h_r_3_49704),
    .O(seg_12_4_sp4_v_b_32_45520)
  );
  LocalMux t5286 (
    .I(seg_12_6_sp4_h_r_7_49708),
    .O(seg_12_6_local_g1_7_49620)
  );
  LocalMux t5287 (
    .I(seg_15_4_sp4_v_b_36_57126),
    .O(seg_15_4_local_g2_4_60870)
  );
  LocalMux t5288 (
    .I(seg_14_7_neigh_op_rgt_2_57350),
    .O(seg_14_7_local_g2_2_57407)
  );
  LocalMux t5289 (
    .I(seg_14_7_neigh_op_rgt_3_57351),
    .O(seg_14_7_local_g3_3_57416)
  );
  CascadeMux t529 (
    .I(net_39254),
    .O(net_39254_cascademuxed)
  );
  LocalMux t5290 (
    .I(seg_14_8_neigh_op_bnr_4_57352),
    .O(seg_14_8_local_g1_4_57524)
  );
  LocalMux t5291 (
    .I(seg_15_7_lutff_6_out_57354),
    .O(seg_15_7_local_g2_6_61241)
  );
  LocalMux t5292 (
    .I(seg_14_9_neigh_op_bnr_2_57473),
    .O(seg_14_9_local_g0_2_57637)
  );
  LocalMux t5293 (
    .I(seg_15_9_neigh_op_bot_2_57473),
    .O(seg_15_9_local_g1_2_61475)
  );
  LocalMux t5294 (
    .I(seg_15_9_neigh_op_bot_3_57474),
    .O(seg_15_9_local_g1_3_61476)
  );
  LocalMux t5295 (
    .I(seg_14_9_neigh_op_bnr_4_57475),
    .O(seg_14_9_local_g0_4_57639)
  );
  LocalMux t5296 (
    .I(seg_15_9_neigh_op_bot_4_57475),
    .O(seg_15_9_local_g0_4_61469)
  );
  LocalMux t5297 (
    .I(seg_2_15_sp4_v_b_19_8656),
    .O(seg_2_15_local_g0_3_13036)
  );
  Span4Mux_v3 t5298 (
    .I(seg_2_12_sp4_h_r_6_12766),
    .O(seg_2_15_sp4_v_b_19_8656)
  );
  Span4Mux_h4 t5299 (
    .I(seg_6_12_sp4_h_r_6_27837),
    .O(seg_2_12_sp4_h_r_6_12766)
  );
  CascadeMux t53 (
    .I(net_9295),
    .O(net_9295_cascademuxed)
  );
  CascadeMux t530 (
    .I(net_39260),
    .O(net_39260_cascademuxed)
  );
  Span4Mux_h4 t5300 (
    .I(seg_10_12_sp4_v_b_1_38587),
    .O(seg_6_12_sp4_h_r_6_27837)
  );
  Span4Mux_v4 t5301 (
    .I(seg_10_8_sp4_h_r_1_42284),
    .O(seg_10_12_sp4_v_b_1_38587)
  );
  Span4Mux_h4 t5302 (
    .I(seg_14_8_sp4_h_r_5_57613),
    .O(seg_10_8_sp4_h_r_1_42284)
  );
  LocalMux t5303 (
    .I(seg_3_8_sp4_h_r_18_12275),
    .O(seg_3_8_local_g1_2_16013)
  );
  Span4Mux_h3 t5304 (
    .I(seg_6_8_sp4_h_r_4_27427),
    .O(seg_3_8_sp4_h_r_18_12275)
  );
  Span4Mux_h4 t5305 (
    .I(seg_10_8_sp4_h_r_1_42284),
    .O(seg_6_8_sp4_h_r_4_27427)
  );
  LocalMux t5306 (
    .I(seg_6_9_sp4_v_b_42_23900),
    .O(seg_6_9_local_g2_2_27467)
  );
  Span4Mux_v1 t5307 (
    .I(seg_6_8_sp4_h_r_1_27422),
    .O(seg_6_9_sp4_v_b_42_23900)
  );
  Span4Mux_h4 t5308 (
    .I(seg_10_8_sp4_h_r_1_42284),
    .O(seg_6_8_sp4_h_r_1_27422)
  );
  LocalMux t5309 (
    .I(seg_6_11_sp4_v_b_18_23900),
    .O(seg_6_11_local_g0_2_27655)
  );
  CascadeMux t531 (
    .I(net_39266),
    .O(net_39266_cascademuxed)
  );
  Span4Mux_v3 t5310 (
    .I(seg_6_8_sp4_h_r_1_27422),
    .O(seg_6_11_sp4_v_b_18_23900)
  );
  LocalMux t5311 (
    .I(seg_6_11_sp4_v_b_20_23902),
    .O(seg_6_11_local_g0_4_27657)
  );
  Span4Mux_v3 t5312 (
    .I(seg_6_8_sp4_h_r_9_27432),
    .O(seg_6_11_sp4_v_b_20_23902)
  );
  Span4Mux_h4 t5313 (
    .I(seg_10_8_sp4_h_r_1_42284),
    .O(seg_6_8_sp4_h_r_9_27432)
  );
  LocalMux t5314 (
    .I(seg_6_12_sp4_h_r_11_27832),
    .O(seg_6_12_local_g1_3_27766)
  );
  Span4Mux_h4 t5315 (
    .I(seg_10_12_sp4_h_r_11_42778),
    .O(seg_6_12_sp4_h_r_11_27832)
  );
  Span4Mux_h4 t5316 (
    .I(seg_14_12_sp4_v_b_11_53921),
    .O(seg_10_12_sp4_h_r_11_42778)
  );
  Span4Mux_v4 t5317 (
    .I(seg_14_8_sp4_h_r_5_57613),
    .O(seg_14_12_sp4_v_b_11_53921)
  );
  LocalMux t5318 (
    .I(seg_13_7_sp4_r_v_b_17_53424),
    .O(seg_13_7_local_g3_1_53584)
  );
  Span4Mux_v1 t5319 (
    .I(seg_14_8_sp4_h_r_11_57609),
    .O(seg_13_7_sp4_r_v_b_17_53424)
  );
  CascadeMux t532 (
    .I(net_39272),
    .O(net_39272_cascademuxed)
  );
  LocalMux t5320 (
    .I(seg_13_7_sp4_v_b_16_49592),
    .O(seg_13_7_local_g1_0_53567)
  );
  Span4Mux_v1 t5321 (
    .I(seg_13_8_sp4_h_r_0_53776),
    .O(seg_13_7_sp4_v_b_16_49592)
  );
  LocalMux t5322 (
    .I(seg_16_11_sp4_r_v_b_23_65413),
    .O(seg_16_11_local_g3_7_65573)
  );
  Span4Mux_v3 t5323 (
    .I(seg_17_8_sp4_h_l_47_53778),
    .O(seg_16_11_sp4_r_v_b_23_65413)
  );
  LocalMux t5324 (
    .I(seg_17_11_sp4_v_b_23_65413),
    .O(seg_17_11_local_g0_7_69380)
  );
  Span4Mux_v3 t5325 (
    .I(seg_17_8_sp4_h_l_47_53778),
    .O(seg_17_11_sp4_v_b_23_65413)
  );
  LocalMux t5326 (
    .I(seg_12_9_sp4_v_b_40_46253),
    .O(seg_12_9_local_g3_0_49998)
  );
  Span4Mux_v1 t5327 (
    .I(seg_12_8_sp4_h_r_5_49952),
    .O(seg_12_9_sp4_v_b_40_46253)
  );
  LocalMux t5328 (
    .I(seg_12_9_sp4_h_r_3_50073),
    .O(seg_12_9_local_g1_3_49985)
  );
  Span4Mux_h4 t5329 (
    .I(seg_16_9_sp4_v_b_10_61213),
    .O(seg_12_9_sp4_h_r_3_50073)
  );
  CascadeMux t533 (
    .I(net_39278),
    .O(net_39278_cascademuxed)
  );
  LocalMux t5330 (
    .I(seg_13_9_sp4_h_r_14_50073),
    .O(seg_13_9_local_g0_6_53811)
  );
  Span4Mux_h3 t5331 (
    .I(seg_16_9_sp4_v_b_10_61213),
    .O(seg_13_9_sp4_h_r_14_50073)
  );
  LocalMux t5332 (
    .I(seg_16_3_sp4_v_b_22_60592),
    .O(seg_16_3_local_g0_6_64564)
  );
  Span4Mux_v1 t5333 (
    .I(seg_16_4_sp4_v_t_38_61081),
    .O(seg_16_3_sp4_v_b_22_60592)
  );
  LocalMux t5334 (
    .I(seg_20_2_sp4_v_b_27_75885),
    .O(seg_20_2_local_g3_3_79155)
  );
  Span4Mux_v2 t5335 (
    .I(seg_20_4_sp4_h_l_38_64780),
    .O(seg_20_2_sp4_v_b_27_75885)
  );
  Span4Mux_h4 t5336 (
    .I(seg_16_4_sp4_v_t_38_61081),
    .O(seg_20_4_sp4_h_l_38_64780)
  );
  LocalMux t5337 (
    .I(seg_20_4_sp4_h_r_6_79476),
    .O(seg_20_4_local_g1_6_79388)
  );
  Span4Mux_h0 t5338 (
    .I(seg_20_4_sp4_h_l_38_64780),
    .O(seg_20_4_sp4_h_r_6_79476)
  );
  LocalMux t5339 (
    .I(seg_15_14_sp4_r_v_b_2_61820),
    .O(seg_15_14_local_g1_2_62090)
  );
  CascadeMux t534 (
    .I(net_39284),
    .O(net_39284_cascademuxed)
  );
  Span4Mux_v4 t5340 (
    .I(seg_16_10_sp4_v_b_11_61335),
    .O(seg_15_14_sp4_r_v_b_2_61820)
  );
  LocalMux t5341 (
    .I(seg_16_11_sp4_v_b_39_61820),
    .O(seg_16_11_local_g2_7_65565)
  );
  Span4Mux_v1 t5342 (
    .I(seg_16_10_sp4_v_b_11_61335),
    .O(seg_16_11_sp4_v_b_39_61820)
  );
  LocalMux t5343 (
    .I(seg_18_2_sp4_h_r_35_64532),
    .O(seg_18_2_local_g2_3_72116)
  );
  Span4Mux_h2 t5344 (
    .I(seg_16_2_sp4_v_t_46_60843),
    .O(seg_18_2_sp4_h_r_35_64532)
  );
  Span4Mux_v4 t5345 (
    .I(seg_16_6_sp4_v_t_46_61335),
    .O(seg_16_2_sp4_v_t_46_60843)
  );
  LocalMux t5346 (
    .I(seg_20_10_sp4_h_r_1_80207),
    .O(seg_20_10_local_g0_1_80113)
  );
  Span4Mux_h0 t5347 (
    .I(seg_20_10_sp4_h_l_40_65520),
    .O(seg_20_10_sp4_h_r_1_80207)
  );
  Span4Mux_h4 t5348 (
    .I(seg_16_10_sp4_v_b_11_61335),
    .O(seg_20_10_sp4_h_l_40_65520)
  );
  LocalMux t5349 (
    .I(seg_6_3_sp4_r_v_b_16_26718),
    .O(seg_6_3_local_g3_0_26861)
  );
  CascadeMux t535 (
    .I(net_39401),
    .O(net_39401_cascademuxed)
  );
  Span4Mux_v1 t5350 (
    .I(seg_7_4_sp4_h_r_0_30298),
    .O(seg_6_3_sp4_r_v_b_16_26718)
  );
  Span4Mux_h4 t5351 (
    .I(seg_11_4_sp4_h_r_0_45622),
    .O(seg_7_4_sp4_h_r_0_30298)
  );
  Span4Mux_h4 t5352 (
    .I(seg_15_4_sp4_v_t_37_57250),
    .O(seg_11_4_sp4_h_r_0_45622)
  );
  LocalMux t5353 (
    .I(seg_6_3_sp4_r_v_b_21_26723),
    .O(seg_6_3_local_g3_5_26866)
  );
  Span4Mux_v1 t5354 (
    .I(seg_7_4_sp4_h_r_3_30303),
    .O(seg_6_3_sp4_r_v_b_21_26723)
  );
  Span4Mux_h4 t5355 (
    .I(seg_11_4_sp4_h_r_0_45622),
    .O(seg_7_4_sp4_h_r_3_30303)
  );
  LocalMux t5356 (
    .I(seg_6_4_sp4_r_v_b_5_26718),
    .O(seg_6_4_local_g1_5_26952)
  );
  Span4Mux_v1 t5357 (
    .I(seg_7_4_sp4_h_r_0_30298),
    .O(seg_6_4_sp4_r_v_b_5_26718)
  );
  LocalMux t5358 (
    .I(seg_2_10_sp4_r_v_b_7_12161),
    .O(seg_2_10_local_g1_7_12433)
  );
  Span4Mux_v1 t5359 (
    .I(seg_3_10_sp4_h_r_7_16352),
    .O(seg_2_10_sp4_r_v_b_7_12161)
  );
  CascadeMux t536 (
    .I(net_39419),
    .O(net_39419_cascademuxed)
  );
  Span4Mux_h4 t5360 (
    .I(seg_7_10_sp4_h_r_4_31042),
    .O(seg_3_10_sp4_h_r_7_16352)
  );
  Span4Mux_h4 t5361 (
    .I(seg_11_10_sp4_h_r_8_46370),
    .O(seg_7_10_sp4_h_r_4_31042)
  );
  Span4Mux_h4 t5362 (
    .I(seg_15_10_sp4_v_b_8_57504),
    .O(seg_11_10_sp4_h_r_8_46370)
  );
  LocalMux t5363 (
    .I(seg_3_14_sp4_v_b_1_12647),
    .O(seg_3_14_local_g0_1_16742)
  );
  Span4Mux_v4 t5364 (
    .I(seg_3_10_sp4_h_r_7_16352),
    .O(seg_3_14_sp4_v_b_1_12647)
  );
  LocalMux t5365 (
    .I(seg_6_9_sp4_r_v_b_12_27331),
    .O(seg_6_9_local_g2_4_27469)
  );
  Span4Mux_v1 t5366 (
    .I(seg_7_10_sp4_h_r_8_31046),
    .O(seg_6_9_sp4_r_v_b_12_27331)
  );
  Span4Mux_h4 t5367 (
    .I(seg_11_10_sp4_h_r_8_46370),
    .O(seg_7_10_sp4_h_r_8_31046)
  );
  LocalMux t5368 (
    .I(seg_6_10_sp4_h_r_42_16352),
    .O(seg_6_10_local_g2_2_27569)
  );
  Span4Mux_h1 t5369 (
    .I(seg_7_10_sp4_h_r_4_31042),
    .O(seg_6_10_sp4_h_r_42_16352)
  );
  CascadeMux t537 (
    .I(net_39506),
    .O(net_39506_cascademuxed)
  );
  LocalMux t5370 (
    .I(seg_17_14_sp4_h_r_34_62176),
    .O(seg_17_14_local_g2_2_69760)
  );
  Span4Mux_h2 t5371 (
    .I(seg_15_14_sp4_v_b_4_57992),
    .O(seg_17_14_sp4_h_r_34_62176)
  );
  Span4Mux_v4 t5372 (
    .I(seg_15_10_sp4_v_b_8_57504),
    .O(seg_15_14_sp4_v_b_4_57992)
  );
  LocalMux t5373 (
    .I(seg_13_7_sp4_h_r_31_46000),
    .O(seg_13_7_local_g3_7_53590)
  );
  Span4Mux_h2 t5374 (
    .I(seg_15_7_sp4_v_t_36_57618),
    .O(seg_13_7_sp4_h_r_31_46000)
  );
  LocalMux t5375 (
    .I(seg_14_11_sp4_r_v_b_1_57618),
    .O(seg_14_11_local_g1_1_57890)
  );
  LocalMux t5376 (
    .I(seg_17_8_sp4_v_b_17_65038),
    .O(seg_17_8_local_g1_1_69013)
  );
  Span4Mux_v1 t5377 (
    .I(seg_17_9_sp4_h_l_41_53905),
    .O(seg_17_8_sp4_v_b_17_65038)
  );
  LocalMux t5378 (
    .I(seg_17_8_sp4_v_b_15_65036),
    .O(seg_17_8_local_g1_7_69019)
  );
  Span4Mux_v1 t5379 (
    .I(seg_17_9_sp4_h_l_45_53909),
    .O(seg_17_8_sp4_v_b_15_65036)
  );
  CascadeMux t538 (
    .I(net_39512),
    .O(net_39512_cascademuxed)
  );
  LocalMux t5380 (
    .I(seg_16_12_sp4_v_b_19_61701),
    .O(seg_16_12_local_g0_3_65668)
  );
  Span4Mux_v3 t5381 (
    .I(seg_16_9_sp4_v_b_3_61204),
    .O(seg_16_12_sp4_v_b_19_61701)
  );
  LocalMux t5382 (
    .I(seg_16_12_sp4_v_b_0_61572),
    .O(seg_16_12_local_g1_0_65673)
  );
  LocalMux t5383 (
    .I(seg_17_8_sp4_h_r_18_65276),
    .O(seg_17_8_local_g0_2_69006)
  );
  Span4Mux_h1 t5384 (
    .I(seg_16_8_sp4_v_t_39_61574),
    .O(seg_17_8_sp4_h_r_18_65276)
  );
  LocalMux t5385 (
    .I(seg_16_12_sp4_v_b_4_61576),
    .O(seg_16_12_local_g1_4_65677)
  );
  LocalMux t5386 (
    .I(seg_15_10_lutff_1_out_57718),
    .O(seg_15_10_local_g1_1_61597)
  );
  LocalMux t5387 (
    .I(seg_15_11_neigh_op_bot_1_57718),
    .O(seg_15_11_local_g1_1_61720)
  );
  LocalMux t5388 (
    .I(seg_15_10_lutff_2_out_57719),
    .O(seg_15_10_local_g3_2_61614)
  );
  LocalMux t5389 (
    .I(seg_15_11_neigh_op_bot_2_57719),
    .O(seg_15_11_local_g0_2_61713)
  );
  CascadeMux t539 (
    .I(net_39518),
    .O(net_39518_cascademuxed)
  );
  LocalMux t5390 (
    .I(seg_15_10_lutff_3_out_57720),
    .O(seg_15_10_local_g2_3_61607)
  );
  LocalMux t5391 (
    .I(seg_15_11_neigh_op_bot_3_57720),
    .O(seg_15_11_local_g0_3_61714)
  );
  LocalMux t5392 (
    .I(seg_15_10_lutff_6_out_57723),
    .O(seg_15_10_local_g1_6_61602)
  );
  LocalMux t5393 (
    .I(seg_15_10_lutff_6_out_57723),
    .O(seg_15_10_local_g2_6_61610)
  );
  LocalMux t5394 (
    .I(seg_15_11_neigh_op_bot_6_57723),
    .O(seg_15_11_local_g1_6_61725)
  );
  LocalMux t5395 (
    .I(seg_15_10_sp4_h_r_26_54026),
    .O(seg_15_10_local_g2_2_61606)
  );
  Span4Mux_h2 t5396 (
    .I(seg_17_10_sp4_h_r_6_69352),
    .O(seg_15_10_sp4_h_r_26_54026)
  );
  Span4Mux_h0 t5397 (
    .I(seg_17_10_sp4_h_l_43_54030),
    .O(seg_17_10_sp4_h_r_6_69352)
  );
  LocalMux t5398 (
    .I(seg_14_12_neigh_op_bnr_0_57840),
    .O(seg_14_12_local_g1_0_58012)
  );
  LocalMux t5399 (
    .I(seg_15_10_neigh_op_top_0_57840),
    .O(seg_15_10_local_g0_0_61588)
  );
  CascadeMux t54 (
    .I(net_9436),
    .O(net_9436_cascademuxed)
  );
  CascadeMux t540 (
    .I(net_39623),
    .O(net_39623_cascademuxed)
  );
  LocalMux t5400 (
    .I(seg_15_10_neigh_op_top_0_57840),
    .O(seg_15_10_local_g1_0_61596)
  );
  LocalMux t5401 (
    .I(seg_15_11_lutff_1_out_57841),
    .O(seg_15_11_local_g3_1_61736)
  );
  LocalMux t5402 (
    .I(seg_15_11_lutff_2_out_57842),
    .O(seg_15_11_local_g3_2_61737)
  );
  LocalMux t5403 (
    .I(seg_16_10_neigh_op_tnl_3_57843),
    .O(seg_16_10_local_g3_3_65446)
  );
  LocalMux t5404 (
    .I(seg_15_11_lutff_4_out_57844),
    .O(seg_15_11_local_g2_4_61731)
  );
  LocalMux t5405 (
    .I(seg_15_12_neigh_op_bot_7_57847),
    .O(seg_15_12_local_g0_7_61841)
  );
  LocalMux t5406 (
    .I(seg_15_14_sp4_v_b_13_58111),
    .O(seg_15_14_local_g1_5_62093)
  );
  Span4Mux_v3 t5407 (
    .I(seg_15_11_sp4_h_r_0_61805),
    .O(seg_15_14_sp4_v_b_13_58111)
  );
  LocalMux t5408 (
    .I(seg_13_14_sp4_r_v_b_22_54290),
    .O(seg_13_14_local_g3_6_54450)
  );
  Span4Mux_v3 t5409 (
    .I(seg_14_11_sp4_h_r_5_57982),
    .O(seg_13_14_sp4_r_v_b_22_54290)
  );
  CascadeMux t541 (
    .I(net_39629),
    .O(net_39629_cascademuxed)
  );
  LocalMux t5410 (
    .I(seg_17_11_sp4_h_r_46_57978),
    .O(seg_17_11_local_g2_6_69395)
  );
  LocalMux t5411 (
    .I(seg_10_11_sp4_h_r_17_38827),
    .O(seg_10_11_local_g1_1_42567)
  );
  Span4Mux_h3 t5412 (
    .I(seg_13_11_sp4_h_r_4_54151),
    .O(seg_10_11_sp4_h_r_17_38827)
  );
  LocalMux t5413 (
    .I(seg_11_11_sp4_r_v_b_0_46127),
    .O(seg_11_11_local_g1_0_46397)
  );
  Span4Mux_v1 t5414 (
    .I(seg_12_11_sp4_h_r_7_50323),
    .O(seg_11_11_sp4_r_v_b_0_46127)
  );
  LocalMux t5415 (
    .I(seg_16_13_sp4_v_b_9_61702),
    .O(seg_16_13_local_g1_1_65797)
  );
  LocalMux t5416 (
    .I(seg_13_14_sp4_h_r_21_50693),
    .O(seg_13_14_local_g1_5_54433)
  );
  Span4Mux_h3 t5417 (
    .I(seg_16_14_sp4_v_b_8_61826),
    .O(seg_13_14_sp4_h_r_21_50693)
  );
  LocalMux t5418 (
    .I(seg_12_12_sp4_h_r_12_46607),
    .O(seg_12_12_local_g1_4_50355)
  );
  Span4Mux_h3 t5419 (
    .I(seg_15_12_sp4_v_b_1_57741),
    .O(seg_12_12_sp4_h_r_12_46607)
  );
  CascadeMux t542 (
    .I(net_39635),
    .O(net_39635_cascademuxed)
  );
  LocalMux t5420 (
    .I(seg_11_14_sp4_h_r_2_46856),
    .O(seg_11_14_local_g1_2_46768)
  );
  Span4Mux_h4 t5421 (
    .I(seg_15_14_sp4_v_b_9_57995),
    .O(seg_11_14_sp4_h_r_2_46856)
  );
  LocalMux t5422 (
    .I(seg_15_12_lutff_1_out_57964),
    .O(seg_15_12_local_g1_1_61843)
  );
  LocalMux t5423 (
    .I(seg_16_13_neigh_op_bnl_2_57965),
    .O(seg_16_13_local_g3_2_65814)
  );
  LocalMux t5424 (
    .I(seg_16_13_neigh_op_bnl_3_57966),
    .O(seg_16_13_local_g2_3_65807)
  );
  LocalMux t5425 (
    .I(seg_16_13_neigh_op_bnl_4_57967),
    .O(seg_16_13_local_g3_4_65816)
  );
  LocalMux t5426 (
    .I(seg_16_11_neigh_op_tnl_6_57969),
    .O(seg_16_11_local_g3_6_65572)
  );
  LocalMux t5427 (
    .I(seg_15_12_lutff_7_out_57970),
    .O(seg_15_12_local_g2_7_61857)
  );
  LocalMux t5428 (
    .I(seg_15_14_sp4_r_v_b_9_61825),
    .O(seg_15_14_local_g2_1_62097)
  );
  LocalMux t5429 (
    .I(seg_18_10_sp4_h_r_42_61691),
    .O(seg_18_10_local_g3_2_73107)
  );
  CascadeMux t543 (
    .I(net_39653),
    .O(net_39653_cascademuxed)
  );
  Span4Mux_h3 t5430 (
    .I(seg_15_10_sp4_v_t_39_57990),
    .O(seg_18_10_sp4_h_r_42_61691)
  );
  LocalMux t5431 (
    .I(seg_15_14_neigh_op_bot_1_58087),
    .O(seg_15_14_local_g0_1_62081)
  );
  LocalMux t5432 (
    .I(seg_15_14_neigh_op_bot_2_58088),
    .O(seg_15_14_local_g0_2_62082)
  );
  LocalMux t5433 (
    .I(seg_15_14_neigh_op_bot_3_58089),
    .O(seg_15_14_local_g0_3_62083)
  );
  LocalMux t5434 (
    .I(seg_15_14_neigh_op_bot_5_58091),
    .O(seg_15_14_local_g0_5_62085)
  );
  LocalMux t5435 (
    .I(seg_15_12_neigh_op_top_7_58093),
    .O(seg_15_12_local_g1_7_61849)
  );
  LocalMux t5436 (
    .I(seg_16_11_sp4_v_b_29_61698),
    .O(seg_16_11_local_g3_5_65571)
  );
  Span4Mux_v2 t5437 (
    .I(seg_16_13_sp4_h_l_40_50567),
    .O(seg_16_11_sp4_v_b_29_61698)
  );
  LocalMux t5438 (
    .I(seg_16_11_sp4_h_r_20_61816),
    .O(seg_16_11_local_g0_4_65546)
  );
  Span4Mux_h1 t5439 (
    .I(seg_15_11_sp4_v_t_41_58115),
    .O(seg_16_11_sp4_h_r_20_61816)
  );
  CascadeMux t544 (
    .I(net_39659),
    .O(net_39659_cascademuxed)
  );
  LocalMux t5440 (
    .I(seg_15_15_neigh_op_bot_1_58210),
    .O(seg_15_15_local_g1_1_62212)
  );
  LocalMux t5441 (
    .I(seg_14_13_neigh_op_tnr_4_58213),
    .O(seg_14_13_local_g2_4_58147)
  );
  LocalMux t5442 (
    .I(seg_15_13_neigh_op_top_5_58214),
    .O(seg_15_13_local_g0_5_61962)
  );
  LocalMux t5443 (
    .I(seg_16_14_sp4_h_r_13_62174),
    .O(seg_16_14_local_g1_5_65924)
  );
  LocalMux t5444 (
    .I(seg_18_31_span4_vert_42_75661),
    .O(seg_18_31_local_g0_2_75679)
  );
  Span4Mux_v1 t5445 (
    .I(seg_18_30_sp4_v_b_11_71457),
    .O(seg_18_31_span4_vert_42_75661)
  );
  Span4Mux_v4 t5446 (
    .I(seg_18_26_sp4_v_b_8_70964),
    .O(seg_18_30_sp4_v_b_11_71457)
  );
  Span4Mux_v4 t5447 (
    .I(seg_18_22_sp4_v_b_0_70464),
    .O(seg_18_26_sp4_v_b_8_70964)
  );
  Span4Mux_v4 t5448 (
    .I(seg_18_18_sp4_v_b_9_69979),
    .O(seg_18_22_sp4_v_b_0_70464)
  );
  Span4Mux_v4 t5449 (
    .I(seg_18_14_sp4_h_l_44_58355),
    .O(seg_18_18_sp4_v_b_9_69979)
  );
  CascadeMux t545 (
    .I(net_39665),
    .O(net_39665_cascademuxed)
  );
  LocalMux t5450 (
    .I(seg_13_31_span4_vert_41_56507),
    .O(seg_13_31_local_g1_1_56533)
  );
  Span4Mux_v1 t5451 (
    .I(seg_13_30_sp4_v_b_1_52294),
    .O(seg_13_31_span4_vert_41_56507)
  );
  Span4Mux_v4 t5452 (
    .I(seg_13_26_sp4_v_b_10_51813),
    .O(seg_13_30_sp4_v_b_1_52294)
  );
  Span4Mux_v4 t5453 (
    .I(seg_13_22_sp4_v_b_2_51313),
    .O(seg_13_26_sp4_v_b_10_51813)
  );
  Span4Mux_v4 t5454 (
    .I(seg_13_18_sp4_v_b_6_50825),
    .O(seg_13_22_sp4_v_b_2_51313)
  );
  Span4Mux_v4 t5455 (
    .I(seg_13_14_sp4_h_r_0_54514),
    .O(seg_13_18_sp4_v_b_6_50825)
  );
  LocalMux t5456 (
    .I(seg_9_0_span4_vert_20_33749),
    .O(seg_9_0_local_g0_4_37403)
  );
  Span4Mux_v2 t5457 (
    .I(seg_9_2_sp4_v_t_43_34025),
    .O(seg_9_0_span4_vert_20_33749)
  );
  Span4Mux_v4 t5458 (
    .I(seg_9_6_sp4_v_t_38_34512),
    .O(seg_9_2_sp4_v_t_43_34025)
  );
  Span4Mux_v4 t5459 (
    .I(seg_9_10_sp4_v_t_37_35003),
    .O(seg_9_6_sp4_v_t_38_34512)
  );
  CascadeMux t546 (
    .I(net_41323),
    .O(net_41323_cascademuxed)
  );
  Span4Mux_v4 t5460 (
    .I(seg_9_14_sp4_h_r_0_39190),
    .O(seg_9_10_sp4_v_t_37_35003)
  );
  Span4Mux_h4 t5461 (
    .I(seg_13_14_sp4_h_r_4_54520),
    .O(seg_9_14_sp4_h_r_0_39190)
  );
  LocalMux t5462 (
    .I(seg_13_31_span4_vert_43_56509),
    .O(seg_13_31_local_g0_3_56527)
  );
  Span4Mux_v1 t5463 (
    .I(seg_13_30_sp4_v_b_10_52305),
    .O(seg_13_31_span4_vert_43_56509)
  );
  Span4Mux_v4 t5464 (
    .I(seg_13_26_sp4_v_b_2_51805),
    .O(seg_13_30_sp4_v_b_10_52305)
  );
  Span4Mux_v4 t5465 (
    .I(seg_13_22_sp4_v_b_6_51317),
    .O(seg_13_26_sp4_v_b_2_51805)
  );
  Span4Mux_v4 t5466 (
    .I(seg_13_18_sp4_v_b_10_50829),
    .O(seg_13_22_sp4_v_b_6_51317)
  );
  Span4Mux_v4 t5467 (
    .I(seg_13_14_sp4_h_r_10_54516),
    .O(seg_13_18_sp4_v_b_10_50829)
  );
  LocalMux t5468 (
    .I(seg_18_14_sp4_h_r_41_62180),
    .O(seg_18_14_local_g2_1_73590)
  );
  LocalMux t5469 (
    .I(seg_16_18_sp4_v_b_11_62319),
    .O(seg_16_18_local_g1_3_66414)
  );
  CascadeMux t547 (
    .I(net_41329),
    .O(net_41329_cascademuxed)
  );
  Span4Mux_v4 t5470 (
    .I(seg_16_14_sp4_h_l_46_50686),
    .O(seg_16_18_sp4_v_b_11_62319)
  );
  LocalMux t5471 (
    .I(seg_15_12_sp4_r_v_b_47_61951),
    .O(seg_15_12_local_g3_7_61865)
  );
  LocalMux t5472 (
    .I(seg_16_13_sp4_h_r_3_65887),
    .O(seg_16_13_local_g1_3_65799)
  );
  Span4Mux_h0 t5473 (
    .I(seg_16_13_sp4_v_t_47_62197),
    .O(seg_16_13_sp4_h_r_3_65887)
  );
  LocalMux t5474 (
    .I(seg_9_0_span4_horz_r_7_33619),
    .O(seg_9_0_local_g0_7_37406)
  );
  IoSpan4Mux t5475 (
    .I(seg_12_0_span4_vert_19_45240),
    .O(seg_9_0_span4_horz_r_7_33619)
  );
  Span4Mux_v2 t5476 (
    .I(seg_12_2_sp4_h_r_1_49208),
    .O(seg_12_0_span4_vert_19_45240)
  );
  Span4Mux_h4 t5477 (
    .I(seg_16_2_sp4_v_t_42_60839),
    .O(seg_12_2_sp4_h_r_1_49208)
  );
  Span4Mux_v4 t5478 (
    .I(seg_16_6_sp4_v_t_42_61331),
    .O(seg_16_2_sp4_v_t_42_60839)
  );
  Span4Mux_v4 t5479 (
    .I(seg_16_10_sp4_v_t_42_61823),
    .O(seg_16_6_sp4_v_t_42_61331)
  );
  CascadeMux t548 (
    .I(net_41365),
    .O(net_41365_cascademuxed)
  );
  LocalMux t5480 (
    .I(seg_15_12_sp4_v_b_34_57998),
    .O(seg_15_12_local_g2_2_61852)
  );
  LocalMux t5481 (
    .I(seg_15_12_sp4_v_b_36_58110),
    .O(seg_15_12_local_g2_4_61854)
  );
  LocalMux t5482 (
    .I(seg_15_15_lutff_1_out_58333),
    .O(seg_15_15_local_g3_1_62228)
  );
  LocalMux t5483 (
    .I(seg_15_15_lutff_2_out_58334),
    .O(seg_15_15_local_g1_2_62213)
  );
  LocalMux t5484 (
    .I(seg_16_14_neigh_op_tnl_3_58335),
    .O(seg_16_14_local_g3_3_65938)
  );
  LocalMux t5485 (
    .I(seg_15_14_neigh_op_top_4_58336),
    .O(seg_15_14_local_g1_4_62092)
  );
  LocalMux t5486 (
    .I(seg_16_13_sp4_v_b_39_62066),
    .O(seg_16_13_local_g3_7_65819)
  );
  LocalMux t5487 (
    .I(seg_9_16_sp4_h_r_18_35614),
    .O(seg_9_16_local_g1_2_39352)
  );
  Span4Mux_h3 t5488 (
    .I(seg_12_16_sp4_h_r_4_50935),
    .O(seg_9_16_sp4_h_r_18_35614)
  );
  Span4Mux_h4 t5489 (
    .I(seg_16_16_sp4_v_b_4_62068),
    .O(seg_12_16_sp4_h_r_4_50935)
  );
  LocalMux t5490 (
    .I(seg_16_13_sp4_v_b_33_61948),
    .O(seg_16_13_local_g3_1_65813)
  );
  LocalMux t5491 (
    .I(seg_15_11_sp4_v_b_20_57749),
    .O(seg_15_11_local_g1_4_61723)
  );
  Span4Mux_v1 t5492 (
    .I(seg_15_12_sp4_v_t_36_58233),
    .O(seg_15_11_sp4_v_b_20_57749)
  );
  LocalMux t5493 (
    .I(seg_10_16_sp4_r_v_b_12_43033),
    .O(seg_10_16_local_g2_4_43193)
  );
  Span4Mux_v1 t5494 (
    .I(seg_11_17_sp4_h_r_1_47222),
    .O(seg_10_16_sp4_r_v_b_12_43033)
  );
  Span4Mux_h4 t5495 (
    .I(seg_15_17_sp4_v_b_8_58365),
    .O(seg_11_17_sp4_h_r_1_47222)
  );
  LocalMux t5496 (
    .I(seg_10_17_sp4_r_v_b_1_43033),
    .O(seg_10_17_local_g1_1_43305)
  );
  Span4Mux_v1 t5497 (
    .I(seg_11_17_sp4_h_r_1_47222),
    .O(seg_10_17_sp4_r_v_b_1_43033)
  );
  LocalMux t5498 (
    .I(seg_11_17_sp4_h_r_1_47222),
    .O(seg_11_17_local_g0_1_47128)
  );
  LocalMux t5499 (
    .I(seg_16_17_neigh_op_bnl_1_58456),
    .O(seg_16_17_local_g2_1_66297)
  );
  CascadeMux t55 (
    .I(net_9625),
    .O(net_9625_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t550 (
    .carryinitin(),
    .carryinitout(t549)
  );
  LocalMux t5500 (
    .I(seg_16_16_neigh_op_lft_2_58457),
    .O(seg_16_16_local_g1_2_66167)
  );
  LocalMux t5501 (
    .I(seg_16_16_neigh_op_lft_4_58459),
    .O(seg_16_16_local_g1_4_66169)
  );
  LocalMux t5502 (
    .I(seg_16_16_neigh_op_lft_5_58460),
    .O(seg_16_16_local_g0_5_66162)
  );
  LocalMux t5503 (
    .I(seg_16_16_neigh_op_lft_7_58462),
    .O(seg_16_16_local_g0_7_66164)
  );
  LocalMux t5504 (
    .I(seg_14_18_sp4_r_v_b_14_58604),
    .O(seg_14_18_local_g2_6_58764)
  );
  LocalMux t5505 (
    .I(seg_14_18_sp4_r_v_b_20_58610),
    .O(seg_14_18_local_g3_4_58770)
  );
  LocalMux t5506 (
    .I(seg_16_17_neigh_op_lft_0_58578),
    .O(seg_16_17_local_g0_0_66280)
  );
  LocalMux t5507 (
    .I(seg_14_16_neigh_op_tnr_2_58580),
    .O(seg_14_16_local_g3_2_58522)
  );
  LocalMux t5508 (
    .I(seg_15_17_lutff_2_out_58580),
    .O(seg_15_17_local_g2_2_62467)
  );
  LocalMux t5509 (
    .I(seg_16_17_neigh_op_lft_4_58582),
    .O(seg_16_17_local_g0_4_66284)
  );
  CascadeMux t551 (
    .I(net_41504),
    .O(net_41504_cascademuxed)
  );
  LocalMux t5510 (
    .I(seg_18_17_sp4_h_r_39_62547),
    .O(seg_18_17_local_g3_7_73973)
  );
  LocalMux t5511 (
    .I(seg_15_15_sp4_v_b_45_58488),
    .O(seg_15_15_local_g3_5_62232)
  );
  LocalMux t5512 (
    .I(seg_15_6_sp4_v_b_11_57013),
    .O(seg_15_6_local_g1_3_61107)
  );
  Span4Mux_v4 t5513 (
    .I(seg_15_2_sp4_h_r_11_60701),
    .O(seg_15_6_sp4_v_b_11_57013)
  );
  LocalMux t5514 (
    .I(seg_16_3_lutff_2_out_60688),
    .O(seg_16_3_local_g1_2_64568)
  );
  LocalMux t5515 (
    .I(seg_4_17_sp12_h_r_0_21031),
    .O(seg_4_17_local_g1_0_20949)
  );
  Span12Mux_h12 t5516 (
    .I(seg_16_17_sp12_v_b_0_64897),
    .O(seg_4_17_sp12_h_r_0_21031)
  );
  Span12Mux_v12 t5517 (
    .I(seg_16_5_sp12_v_b_0_64260),
    .O(seg_16_17_sp12_v_b_0_64897)
  );
  LocalMux t5518 (
    .I(seg_4_7_sp4_r_v_b_10_19459),
    .O(seg_4_7_local_g2_2_19729)
  );
  Span4Mux_v4 t5519 (
    .I(seg_5_3_sp4_h_r_4_23150),
    .O(seg_4_7_sp4_r_v_b_10_19459)
  );
  Span4Mux_h4 t5520 (
    .I(seg_9_3_sp4_h_r_1_37838),
    .O(seg_5_3_sp4_h_r_4_23150)
  );
  Span4Mux_h4 t5521 (
    .I(seg_13_3_sp4_h_r_1_53162),
    .O(seg_9_3_sp4_h_r_1_37838)
  );
  LocalMux t5522 (
    .I(seg_4_18_sp4_r_v_b_19_20931),
    .O(seg_4_18_local_g3_3_21091)
  );
  Span4Mux_v3 t5523 (
    .I(seg_5_15_sp4_h_r_0_24620),
    .O(seg_4_18_sp4_r_v_b_19_20931)
  );
  Span4Mux_h4 t5524 (
    .I(seg_9_15_sp4_h_r_4_39319),
    .O(seg_5_15_sp4_h_r_0_24620)
  );
  Span4Mux_h4 t5525 (
    .I(seg_13_15_sp4_v_b_4_50454),
    .O(seg_9_15_sp4_h_r_4_39319)
  );
  Span4Mux_v4 t5526 (
    .I(seg_13_11_sp4_v_b_1_49957),
    .O(seg_13_15_sp4_v_b_4_50454)
  );
  Span4Mux_v4 t5527 (
    .I(seg_13_7_sp4_v_b_1_49465),
    .O(seg_13_11_sp4_v_b_1_49957)
  );
  Span4Mux_v4 t5528 (
    .I(seg_13_3_sp4_h_r_1_53162),
    .O(seg_13_7_sp4_v_b_1_49465)
  );
  LocalMux t5529 (
    .I(seg_10_19_sp4_h_r_18_39814),
    .O(seg_10_19_local_g0_2_43544)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t553 (
    .carryinitin(),
    .carryinitout(t552)
  );
  Span4Mux_h3 t5530 (
    .I(seg_13_19_sp4_v_b_7_50947),
    .O(seg_10_19_sp4_h_r_18_39814)
  );
  Span4Mux_v4 t5531 (
    .I(seg_13_15_sp4_v_b_4_50454),
    .O(seg_13_19_sp4_v_b_7_50947)
  );
  LocalMux t5532 (
    .I(seg_20_7_sp4_v_b_10_76206),
    .O(seg_20_7_local_g0_2_79745)
  );
  Span4Mux_v4 t5533 (
    .I(seg_20_3_sp4_h_r_4_79351),
    .O(seg_20_7_sp4_v_b_10_76206)
  );
  Span4Mux_h0 t5534 (
    .I(seg_20_3_sp4_h_l_41_64658),
    .O(seg_20_3_sp4_h_r_4_79351)
  );
  LocalMux t5535 (
    .I(seg_16_11_sp4_v_b_2_61451),
    .O(seg_16_11_local_g0_2_65544)
  );
  Span4Mux_v4 t5536 (
    .I(seg_16_7_sp4_v_b_6_60963),
    .O(seg_16_11_sp4_v_b_2_61451)
  );
  Span4Mux_v4 t5537 (
    .I(seg_16_3_sp4_h_r_6_64660),
    .O(seg_16_7_sp4_v_b_6_60963)
  );
  LocalMux t5538 (
    .I(seg_20_4_sp4_v_b_43_76202),
    .O(seg_20_4_local_g3_3_79401)
  );
  Span4Mux_v1 t5539 (
    .I(seg_20_3_sp4_h_l_43_64660),
    .O(seg_20_4_sp4_v_b_43_76202)
  );
  CascadeMux t554 (
    .I(net_41615),
    .O(net_41615_cascademuxed)
  );
  LocalMux t5540 (
    .I(seg_20_10_sp4_v_b_18_76609),
    .O(seg_20_10_local_g0_2_80114)
  );
  Span4Mux_v3 t5541 (
    .I(seg_20_7_sp4_v_b_11_76205),
    .O(seg_20_10_sp4_v_b_18_76609)
  );
  Span4Mux_v4 t5542 (
    .I(seg_20_3_sp4_h_l_43_64660),
    .O(seg_20_7_sp4_v_b_11_76205)
  );
  LocalMux t5543 (
    .I(seg_17_11_sp4_v_b_19_65409),
    .O(seg_17_11_local_g1_3_69384)
  );
  Span4Mux_v3 t5544 (
    .I(seg_17_8_sp4_v_b_10_64921),
    .O(seg_17_11_sp4_v_b_19_65409)
  );
  Span4Mux_v4 t5545 (
    .I(seg_17_4_sp4_v_b_10_64424),
    .O(seg_17_8_sp4_v_b_10_64921)
  );
  LocalMux t5546 (
    .I(seg_20_6_sp4_h_r_43_68860),
    .O(seg_20_6_local_g3_3_79647)
  );
  Span4Mux_h3 t5547 (
    .I(seg_17_6_sp4_v_b_0_64665),
    .O(seg_20_6_sp4_h_r_43_68860)
  );
  LocalMux t5548 (
    .I(seg_5_16_sp4_h_r_18_20921),
    .O(seg_5_16_local_g0_2_24651)
  );
  Span4Mux_h3 t5549 (
    .I(seg_8_16_sp4_h_r_4_35611),
    .O(seg_5_16_sp4_h_r_18_20921)
  );
  CascadeMux t555 (
    .I(net_41627),
    .O(net_41627_cascademuxed)
  );
  Span4Mux_h4 t5550 (
    .I(seg_12_16_sp4_v_b_4_46746),
    .O(seg_8_16_sp4_h_r_4_35611)
  );
  Span4Mux_v4 t5551 (
    .I(seg_12_12_sp4_h_r_10_50439),
    .O(seg_12_16_sp4_v_b_4_46746)
  );
  Span4Mux_h4 t5552 (
    .I(seg_16_12_sp4_v_b_5_61575),
    .O(seg_12_12_sp4_h_r_10_50439)
  );
  Span4Mux_v4 t5553 (
    .I(seg_16_8_sp4_v_b_5_61083),
    .O(seg_16_12_sp4_v_b_5_61575)
  );
  Span4Mux_v4 t5554 (
    .I(seg_16_4_sp4_v_b_9_60590),
    .O(seg_16_8_sp4_v_b_5_61083)
  );
  LocalMux t5555 (
    .I(seg_7_15_sp4_r_v_b_19_31424),
    .O(seg_7_15_local_g3_3_31584)
  );
  Span4Mux_v3 t5556 (
    .I(seg_8_12_sp4_h_r_6_35121),
    .O(seg_7_15_sp4_r_v_b_19_31424)
  );
  Span4Mux_h4 t5557 (
    .I(seg_12_12_sp4_h_r_10_50439),
    .O(seg_8_12_sp4_h_r_6_35121)
  );
  LocalMux t5558 (
    .I(seg_8_16_sp4_h_r_3_35610),
    .O(seg_8_16_local_g1_3_35522)
  );
  Span4Mux_h4 t5559 (
    .I(seg_12_16_sp4_v_b_10_46752),
    .O(seg_8_16_sp4_h_r_3_35610)
  );
  CascadeMux t556 (
    .I(net_41633),
    .O(net_41633_cascademuxed)
  );
  Span4Mux_v4 t5560 (
    .I(seg_12_12_sp4_h_r_10_50439),
    .O(seg_12_16_sp4_v_b_10_46752)
  );
  LocalMux t5561 (
    .I(seg_3_18_sp4_r_v_b_3_16972),
    .O(seg_3_18_local_g1_3_17244)
  );
  Span4Mux_v4 t5562 (
    .I(seg_4_14_sp4_h_r_9_20677),
    .O(seg_3_18_sp4_r_v_b_3_16972)
  );
  Span4Mux_h4 t5563 (
    .I(seg_8_14_sp4_h_r_6_35367),
    .O(seg_4_14_sp4_h_r_9_20677)
  );
  Span4Mux_h4 t5564 (
    .I(seg_12_14_sp4_v_b_6_46502),
    .O(seg_8_14_sp4_h_r_6_35367)
  );
  Span4Mux_v4 t5565 (
    .I(seg_12_10_sp4_v_b_6_46010),
    .O(seg_12_14_sp4_v_b_6_46502)
  );
  Span4Mux_v4 t5566 (
    .I(seg_12_6_sp4_h_r_6_49707),
    .O(seg_12_10_sp4_v_b_6_46010)
  );
  Span4Mux_h4 t5567 (
    .I(seg_16_6_sp4_v_b_1_60833),
    .O(seg_12_6_sp4_h_r_6_49707)
  );
  LocalMux t5568 (
    .I(seg_15_6_sp4_h_r_43_49707),
    .O(seg_15_6_local_g3_3_61123)
  );
  Span4Mux_h1 t5569 (
    .I(seg_16_6_sp4_v_b_1_60833),
    .O(seg_15_6_sp4_h_r_43_49707)
  );
  CascadeMux t557 (
    .I(net_41645),
    .O(net_41645_cascademuxed)
  );
  LocalMux t5570 (
    .I(seg_15_18_sp4_r_v_b_3_62311),
    .O(seg_15_18_local_g1_3_62583)
  );
  Span4Mux_v4 t5571 (
    .I(seg_16_14_sp4_v_b_0_61818),
    .O(seg_15_18_sp4_r_v_b_3_62311)
  );
  Span4Mux_v4 t5572 (
    .I(seg_16_10_sp4_v_b_9_61333),
    .O(seg_16_14_sp4_v_b_0_61818)
  );
  Span4Mux_v4 t5573 (
    .I(seg_16_6_sp4_v_b_1_60833),
    .O(seg_16_10_sp4_v_b_9_61333)
  );
  LocalMux t5574 (
    .I(seg_15_14_sp4_r_v_b_3_61819),
    .O(seg_15_14_local_g1_3_62091)
  );
  Span4Mux_v4 t5575 (
    .I(seg_16_10_sp4_v_b_3_61327),
    .O(seg_15_14_sp4_r_v_b_3_61819)
  );
  Span4Mux_v4 t5576 (
    .I(seg_16_6_sp4_v_b_3_60835),
    .O(seg_16_10_sp4_v_b_3_61327)
  );
  LocalMux t5577 (
    .I(seg_16_6_sp4_r_v_b_3_64666),
    .O(seg_16_6_local_g1_3_64938)
  );
  LocalMux t5578 (
    .I(seg_16_6_sp4_r_v_b_11_64674),
    .O(seg_16_6_local_g2_3_64946)
  );
  LocalMux t5579 (
    .I(seg_16_6_sp4_r_v_b_17_64792),
    .O(seg_16_6_local_g3_1_64952)
  );
  LocalMux t5580 (
    .I(seg_16_6_sp4_r_v_b_21_64796),
    .O(seg_16_6_local_g3_5_64956)
  );
  LocalMux t5581 (
    .I(seg_16_6_sp4_v_b_12_60956),
    .O(seg_16_6_local_g0_4_64931)
  );
  LocalMux t5582 (
    .I(seg_16_6_sp4_v_b_14_60958),
    .O(seg_16_6_local_g0_6_64933)
  );
  LocalMux t5583 (
    .I(seg_16_6_sp4_v_b_22_60966),
    .O(seg_16_6_local_g1_6_64941)
  );
  LocalMux t5584 (
    .I(seg_16_4_neigh_op_top_4_60936),
    .O(seg_16_4_local_g0_4_64685)
  );
  LocalMux t5585 (
    .I(seg_16_6_neigh_op_bot_5_60937),
    .O(seg_16_6_local_g0_5_64932)
  );
  LocalMux t5586 (
    .I(seg_16_4_neigh_op_top_6_60938),
    .O(seg_16_4_local_g1_6_64695)
  );
  LocalMux t5587 (
    .I(seg_16_4_neigh_op_top_7_60939),
    .O(seg_16_4_local_g1_7_64696)
  );
  LocalMux t5588 (
    .I(seg_16_7_sp4_r_v_b_15_64913),
    .O(seg_16_7_local_g2_7_65073)
  );
  LocalMux t5589 (
    .I(seg_16_7_sp4_v_b_8_60965),
    .O(seg_16_7_local_g0_0_65050)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t559 (
    .carryinitin(),
    .carryinitout(t558)
  );
  LocalMux t5590 (
    .I(seg_16_7_sp4_v_b_10_60967),
    .O(seg_16_7_local_g0_2_65052)
  );
  LocalMux t5591 (
    .I(seg_16_7_sp4_v_b_12_61079),
    .O(seg_16_7_local_g1_4_65062)
  );
  LocalMux t5592 (
    .I(seg_16_8_sp4_v_b_7_61085),
    .O(seg_16_8_local_g0_7_65180)
  );
  LocalMux t5593 (
    .I(seg_14_8_sp4_r_v_b_27_57497),
    .O(seg_14_8_local_g1_3_57523)
  );
  Span4Mux_v2 t5594 (
    .I(seg_15_6_sp4_h_r_9_61201),
    .O(seg_14_8_sp4_r_v_b_27_57497)
  );
  LocalMux t5595 (
    .I(seg_10_10_sp4_v_b_2_38344),
    .O(seg_10_10_local_g1_2_42445)
  );
  Span4Mux_v4 t5596 (
    .I(seg_10_6_sp4_h_r_8_42047),
    .O(seg_10_10_sp4_v_b_2_38344)
  );
  Span4Mux_h4 t5597 (
    .I(seg_14_6_sp4_h_r_0_57360),
    .O(seg_10_6_sp4_h_r_8_42047)
  );
  LocalMux t5598 (
    .I(seg_14_8_sp4_v_b_34_53676),
    .O(seg_14_8_local_g3_2_57538)
  );
  Span4Mux_v2 t5599 (
    .I(seg_14_6_sp4_h_r_4_57366),
    .O(seg_14_8_sp4_v_b_34_53676)
  );
  CascadeMux t56 (
    .I(net_9748),
    .O(net_9748_cascademuxed)
  );
  CascadeMux t560 (
    .I(net_41732),
    .O(net_41732_cascademuxed)
  );
  LocalMux t5600 (
    .I(seg_14_7_sp4_h_r_23_53655),
    .O(seg_14_7_local_g1_7_57404)
  );
  Span4Mux_h3 t5601 (
    .I(seg_17_7_sp4_v_b_10_64798),
    .O(seg_14_7_sp4_h_r_23_53655)
  );
  LocalMux t5602 (
    .I(seg_14_8_sp4_h_r_17_53782),
    .O(seg_14_8_local_g0_1_57513)
  );
  Span4Mux_h3 t5603 (
    .I(seg_17_8_sp4_v_b_11_64920),
    .O(seg_14_8_sp4_h_r_17_53782)
  );
  LocalMux t5604 (
    .I(seg_16_9_sp4_v_b_7_61208),
    .O(seg_16_9_local_g0_7_65303)
  );
  LocalMux t5605 (
    .I(seg_14_13_sp4_h_r_26_50564),
    .O(seg_14_13_local_g2_2_58145)
  );
  Span4Mux_h2 t5606 (
    .I(seg_16_13_sp4_v_b_2_61697),
    .O(seg_14_13_sp4_h_r_26_50564)
  );
  Span4Mux_v4 t5607 (
    .I(seg_16_9_sp4_v_b_11_61212),
    .O(seg_16_13_sp4_v_b_2_61697)
  );
  LocalMux t5608 (
    .I(seg_16_7_lutff_3_out_61181),
    .O(seg_16_7_local_g0_3_65053)
  );
  LocalMux t5609 (
    .I(seg_16_7_lutff_4_out_61182),
    .O(seg_16_7_local_g2_4_65070)
  );
  CascadeMux t561 (
    .I(net_41750),
    .O(net_41750_cascademuxed)
  );
  LocalMux t5610 (
    .I(seg_15_15_sp4_r_v_b_3_61942),
    .O(seg_15_15_local_g1_3_62214)
  );
  Span4Mux_v4 t5611 (
    .I(seg_16_11_sp4_v_b_0_61449),
    .O(seg_15_15_sp4_r_v_b_3_61942)
  );
  Span4Mux_v4 t5612 (
    .I(seg_16_7_sp4_h_r_0_65144),
    .O(seg_16_11_sp4_v_b_0_61449)
  );
  LocalMux t5613 (
    .I(seg_12_10_sp4_v_b_21_46135),
    .O(seg_12_10_local_g1_5_50110)
  );
  Span4Mux_v3 t5614 (
    .I(seg_12_7_sp4_h_r_2_49826),
    .O(seg_12_10_sp4_v_b_21_46135)
  );
  Span4Mux_h4 t5615 (
    .I(seg_16_7_sp4_h_r_2_65148),
    .O(seg_12_7_sp4_h_r_2_49826)
  );
  LocalMux t5616 (
    .I(seg_14_13_sp4_r_v_b_33_58118),
    .O(seg_14_13_local_g2_1_58144)
  );
  Span4Mux_v2 t5617 (
    .I(seg_15_11_sp4_v_b_9_57626),
    .O(seg_14_13_sp4_r_v_b_33_58118)
  );
  Span4Mux_v4 t5618 (
    .I(seg_15_7_sp4_h_r_9_61324),
    .O(seg_15_11_sp4_v_b_9_57626)
  );
  LocalMux t5619 (
    .I(seg_18_7_sp4_h_r_46_61316),
    .O(seg_18_7_local_g2_6_72734)
  );
  CascadeMux t562 (
    .I(net_41774),
    .O(net_41774_cascademuxed)
  );
  LocalMux t5620 (
    .I(seg_18_7_sp4_h_r_6_72814),
    .O(seg_18_7_local_g0_6_72718)
  );
  Span4Mux_h0 t5621 (
    .I(seg_18_7_sp4_h_l_43_57491),
    .O(seg_18_7_sp4_h_r_6_72814)
  );
  LocalMux t5622 (
    .I(seg_10_16_sp4_h_r_22_39439),
    .O(seg_10_16_local_g1_6_43187)
  );
  Span4Mux_h3 t5623 (
    .I(seg_13_16_sp4_h_r_8_54770),
    .O(seg_10_16_sp4_h_r_22_39439)
  );
  Span4Mux_h4 t5624 (
    .I(seg_17_16_sp4_v_b_3_65896),
    .O(seg_13_16_sp4_h_r_8_54770)
  );
  Span4Mux_v4 t5625 (
    .I(seg_17_12_sp4_v_b_3_65404),
    .O(seg_17_16_sp4_v_b_3_65896)
  );
  Span4Mux_v4 t5626 (
    .I(seg_17_8_sp4_v_b_0_64911),
    .O(seg_17_12_sp4_v_b_3_65404)
  );
  LocalMux t5627 (
    .I(seg_10_17_sp4_h_r_22_39562),
    .O(seg_10_17_local_g0_6_43302)
  );
  Span4Mux_h3 t5628 (
    .I(seg_13_17_sp4_h_r_11_54886),
    .O(seg_10_17_sp4_h_r_22_39562)
  );
  Span4Mux_h4 t5629 (
    .I(seg_17_17_sp4_v_b_11_66027),
    .O(seg_13_17_sp4_h_r_11_54886)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t563 (
    .carryinitin(net_45602),
    .carryinitout(net_45646)
  );
  Span4Mux_v4 t5630 (
    .I(seg_17_13_sp4_v_b_8_65534),
    .O(seg_17_17_sp4_v_b_11_66027)
  );
  Span4Mux_v4 t5631 (
    .I(seg_17_9_sp4_v_b_5_65037),
    .O(seg_17_13_sp4_v_b_8_65534)
  );
  LocalMux t5632 (
    .I(seg_9_16_sp4_v_b_34_35505),
    .O(seg_9_16_local_g2_2_39360)
  );
  Span4Mux_v2 t5633 (
    .I(seg_9_14_sp4_v_b_2_35005),
    .O(seg_9_16_sp4_v_b_34_35505)
  );
  Span4Mux_v4 t5634 (
    .I(seg_9_10_sp4_h_r_8_38708),
    .O(seg_9_14_sp4_v_b_2_35005)
  );
  Span4Mux_h4 t5635 (
    .I(seg_13_10_sp4_h_r_8_54032),
    .O(seg_9_10_sp4_h_r_8_38708)
  );
  Span4Mux_h4 t5636 (
    .I(seg_17_10_sp4_v_b_8_65165),
    .O(seg_13_10_sp4_h_r_8_54032)
  );
  LocalMux t5637 (
    .I(seg_9_17_sp4_v_b_23_35505),
    .O(seg_9_17_local_g1_7_39480)
  );
  Span4Mux_v3 t5638 (
    .I(seg_9_14_sp4_v_b_2_35005),
    .O(seg_9_17_sp4_v_b_23_35505)
  );
  LocalMux t5639 (
    .I(seg_11_8_sp4_r_v_b_15_45883),
    .O(seg_11_8_local_g2_7_46043)
  );
  CascadeMux t564 (
    .I(net_42107),
    .O(net_42107_cascademuxed)
  );
  Span4Mux_v1 t5640 (
    .I(seg_12_9_sp4_h_r_2_50072),
    .O(seg_11_8_sp4_r_v_b_15_45883)
  );
  Span4Mux_h4 t5641 (
    .I(seg_16_9_sp4_v_b_2_61205),
    .O(seg_12_9_sp4_h_r_2_50072)
  );
  LocalMux t5642 (
    .I(seg_15_8_neigh_op_rgt_0_61301),
    .O(seg_15_8_local_g3_0_61366)
  );
  LocalMux t5643 (
    .I(seg_12_10_sp4_h_r_3_50196),
    .O(seg_12_10_local_g0_3_50100)
  );
  Span4Mux_h4 t5644 (
    .I(seg_16_10_sp4_v_b_10_61336),
    .O(seg_12_10_sp4_h_r_3_50196)
  );
  LocalMux t5645 (
    .I(seg_15_11_sp4_r_v_b_5_61452),
    .O(seg_15_11_local_g1_5_61724)
  );
  LocalMux t5646 (
    .I(seg_15_9_neigh_op_rgt_4_61428),
    .O(seg_15_9_local_g2_4_61485)
  );
  LocalMux t5647 (
    .I(seg_15_9_neigh_op_rgt_7_61431),
    .O(seg_15_9_local_g3_7_61496)
  );
  LocalMux t5648 (
    .I(seg_11_9_sp12_h_r_3_42402),
    .O(seg_11_9_local_g1_3_46154)
  );
  LocalMux t5649 (
    .I(seg_13_10_sp4_r_v_b_37_54035),
    .O(seg_13_10_local_g2_5_53949)
  );
  CascadeMux t565 (
    .I(net_42125),
    .O(net_42125_cascademuxed)
  );
  Span4Mux_v1 t5650 (
    .I(seg_14_9_sp4_h_r_0_57729),
    .O(seg_13_10_sp4_r_v_b_37_54035)
  );
  LocalMux t5651 (
    .I(seg_13_12_sp4_r_v_b_13_54035),
    .O(seg_13_12_local_g2_5_54195)
  );
  Span4Mux_v3 t5652 (
    .I(seg_14_9_sp4_h_r_0_57729),
    .O(seg_13_12_sp4_r_v_b_13_54035)
  );
  LocalMux t5653 (
    .I(seg_13_12_sp4_r_v_b_17_54039),
    .O(seg_13_12_local_g3_1_54199)
  );
  Span4Mux_v3 t5654 (
    .I(seg_14_9_sp4_h_r_10_57731),
    .O(seg_13_12_sp4_r_v_b_17_54039)
  );
  LocalMux t5655 (
    .I(seg_13_13_sp4_r_v_b_4_54039),
    .O(seg_13_13_local_g1_4_54309)
  );
  Span4Mux_v4 t5656 (
    .I(seg_14_9_sp4_h_r_10_57731),
    .O(seg_13_13_sp4_r_v_b_4_54039)
  );
  LocalMux t5657 (
    .I(seg_12_11_sp4_r_v_b_31_50209),
    .O(seg_12_11_local_g1_7_50235)
  );
  Span4Mux_v2 t5658 (
    .I(seg_13_9_sp4_h_r_7_53908),
    .O(seg_12_11_sp4_r_v_b_31_50209)
  );
  LocalMux t5659 (
    .I(seg_13_11_sp4_v_b_31_50209),
    .O(seg_13_11_local_g3_7_54082)
  );
  CascadeMux t566 (
    .I(net_42248),
    .O(net_42248_cascademuxed)
  );
  Span4Mux_v2 t5660 (
    .I(seg_13_9_sp4_h_r_7_53908),
    .O(seg_13_11_sp4_v_b_31_50209)
  );
  LocalMux t5661 (
    .I(seg_13_13_sp4_v_b_7_50209),
    .O(seg_13_13_local_g0_7_54304)
  );
  Span4Mux_v4 t5662 (
    .I(seg_13_9_sp4_h_r_7_53908),
    .O(seg_13_13_sp4_v_b_7_50209)
  );
  LocalMux t5663 (
    .I(seg_12_9_sp4_r_v_b_11_49721),
    .O(seg_12_9_local_g2_3_49993)
  );
  Span4Mux_v1 t5664 (
    .I(seg_13_9_sp4_h_r_11_53902),
    .O(seg_12_9_sp4_r_v_b_11_49721)
  );
  LocalMux t5665 (
    .I(seg_13_7_sp4_v_b_35_49721),
    .O(seg_13_7_local_g2_3_53578)
  );
  Span4Mux_v2 t5666 (
    .I(seg_13_9_sp4_h_r_11_53902),
    .O(seg_13_7_sp4_v_b_35_49721)
  );
  LocalMux t5667 (
    .I(seg_13_9_sp4_h_r_11_53902),
    .O(seg_13_9_local_g1_3_53816)
  );
  LocalMux t5668 (
    .I(seg_14_11_sp4_h_r_19_54153),
    .O(seg_14_11_local_g0_3_57884)
  );
  Span4Mux_h3 t5669 (
    .I(seg_17_11_sp4_v_b_1_65279),
    .O(seg_14_11_sp4_h_r_19_54153)
  );
  CascadeMux t567 (
    .I(net_42365),
    .O(net_42365_cascademuxed)
  );
  LocalMux t5670 (
    .I(seg_16_5_sp4_v_b_17_60838),
    .O(seg_16_5_local_g0_1_64805)
  );
  Span4Mux_v1 t5671 (
    .I(seg_16_6_sp4_v_t_36_61325),
    .O(seg_16_5_sp4_v_b_17_60838)
  );
  LocalMux t5672 (
    .I(seg_12_11_sp4_h_r_10_50316),
    .O(seg_12_11_local_g0_2_50222)
  );
  Span4Mux_h4 t5673 (
    .I(seg_16_11_sp4_v_b_10_61459),
    .O(seg_12_11_sp4_h_r_10_50316)
  );
  LocalMux t5674 (
    .I(seg_13_11_sp4_h_r_23_50316),
    .O(seg_13_11_local_g0_7_54058)
  );
  Span4Mux_h3 t5675 (
    .I(seg_16_11_sp4_v_b_10_61459),
    .O(seg_13_11_sp4_h_r_23_50316)
  );
  LocalMux t5676 (
    .I(seg_13_12_sp4_h_r_13_50437),
    .O(seg_13_12_local_g0_5_54179)
  );
  Span4Mux_h3 t5677 (
    .I(seg_16_12_sp4_v_b_7_61577),
    .O(seg_13_12_sp4_h_r_13_50437)
  );
  LocalMux t5678 (
    .I(seg_16_11_neigh_op_bot_1_61548),
    .O(seg_16_11_local_g0_1_65543)
  );
  LocalMux t5679 (
    .I(seg_25_11_sp4_h_r_0_100236),
    .O(seg_25_11_local_g0_0_100150)
  );
  CascadeMux t568 (
    .I(net_42470),
    .O(net_42470_cascademuxed)
  );
  Span4Mux_h0 t5680 (
    .I(seg_25_11_sp4_h_l_41_84166),
    .O(seg_25_11_sp4_h_r_0_100236)
  );
  Span4Mux_h4 t5681 (
    .I(seg_21_11_sp4_h_l_41_69473),
    .O(seg_25_11_sp4_h_l_41_84166)
  );
  Span4Mux_h4 t5682 (
    .I(seg_17_11_sp4_v_b_4_65284),
    .O(seg_21_11_sp4_h_l_41_69473)
  );
  LocalMux t5683 (
    .I(seg_25_11_sp4_h_r_4_100242),
    .O(seg_25_11_local_g0_4_100154)
  );
  Span4Mux_h0 t5684 (
    .I(seg_25_11_sp4_h_l_45_84170),
    .O(seg_25_11_sp4_h_r_4_100242)
  );
  Span4Mux_h4 t5685 (
    .I(seg_21_11_sp4_h_l_45_69477),
    .O(seg_25_11_sp4_h_l_45_84170)
  );
  Span4Mux_h4 t5686 (
    .I(seg_17_11_sp4_v_b_8_65288),
    .O(seg_21_11_sp4_h_l_45_69477)
  );
  LocalMux t5687 (
    .I(seg_25_12_sp4_v_b_36_95952),
    .O(seg_25_12_local_g2_4_100320)
  );
  Span4Mux_v1 t5688 (
    .I(seg_25_11_sp4_h_l_45_84170),
    .O(seg_25_12_sp4_v_b_36_95952)
  );
  LocalMux t5689 (
    .I(seg_25_11_sp4_h_r_6_100244),
    .O(seg_25_11_local_g0_6_100156)
  );
  CascadeMux t569 (
    .I(net_42500),
    .O(net_42500_cascademuxed)
  );
  Span4Mux_h0 t5690 (
    .I(seg_25_11_sp4_h_l_43_84168),
    .O(seg_25_11_sp4_h_r_6_100244)
  );
  Span4Mux_h4 t5691 (
    .I(seg_21_11_sp4_h_l_47_69469),
    .O(seg_25_11_sp4_h_l_43_84168)
  );
  Span4Mux_h4 t5692 (
    .I(seg_17_11_sp4_v_b_10_65290),
    .O(seg_21_11_sp4_h_l_47_69469)
  );
  LocalMux t5693 (
    .I(seg_25_11_sp4_v_b_21_95544),
    .O(seg_25_11_local_g0_5_100155)
  );
  Span4Mux_v1 t5694 (
    .I(seg_25_12_sp4_h_l_45_84293),
    .O(seg_25_11_sp4_v_b_21_95544)
  );
  Span4Mux_h4 t5695 (
    .I(seg_21_12_sp4_h_l_40_69597),
    .O(seg_25_12_sp4_h_l_45_84293)
  );
  Span4Mux_h4 t5696 (
    .I(seg_17_12_sp4_v_b_5_65406),
    .O(seg_21_12_sp4_h_l_40_69597)
  );
  LocalMux t5697 (
    .I(seg_25_12_sp4_h_r_4_100393),
    .O(seg_25_12_local_g1_4_100312)
  );
  Span4Mux_h0 t5698 (
    .I(seg_25_12_sp4_h_l_45_84293),
    .O(seg_25_12_sp4_h_r_4_100393)
  );
  LocalMux t5699 (
    .I(seg_25_11_sp4_v_b_14_95537),
    .O(seg_25_11_local_g1_6_100164)
  );
  CascadeMux t57 (
    .I(net_9913),
    .O(net_9913_cascademuxed)
  );
  CascadeMux t570 (
    .I(net_42506),
    .O(net_42506_cascademuxed)
  );
  Span4Mux_v1 t5700 (
    .I(seg_25_12_sp4_h_l_38_84288),
    .O(seg_25_11_sp4_v_b_14_95537)
  );
  Span4Mux_h4 t5701 (
    .I(seg_21_12_sp4_h_l_42_69599),
    .O(seg_25_12_sp4_h_l_38_84288)
  );
  Span4Mux_h4 t5702 (
    .I(seg_17_12_sp4_v_b_7_65408),
    .O(seg_21_12_sp4_h_l_42_69599)
  );
  LocalMux t5703 (
    .I(seg_25_12_sp4_h_r_3_100392),
    .O(seg_25_12_local_g0_3_100303)
  );
  Span4Mux_h0 t5704 (
    .I(seg_25_12_sp4_h_l_38_84288),
    .O(seg_25_12_sp4_h_r_3_100392)
  );
  LocalMux t5705 (
    .I(seg_25_12_sp4_h_r_2_100391),
    .O(seg_25_12_local_g0_2_100302)
  );
  Span4Mux_h0 t5706 (
    .I(seg_25_12_sp4_h_l_46_84286),
    .O(seg_25_12_sp4_h_r_2_100391)
  );
  Span4Mux_h4 t5707 (
    .I(seg_21_12_sp4_h_l_38_69595),
    .O(seg_25_12_sp4_h_l_46_84286)
  );
  Span4Mux_h4 t5708 (
    .I(seg_17_12_sp4_v_b_9_65410),
    .O(seg_21_12_sp4_h_l_38_69595)
  );
  LocalMux t5709 (
    .I(seg_25_12_sp4_v_b_21_95683),
    .O(seg_25_12_local_g1_5_100313)
  );
  CascadeMux t571 (
    .I(net_42512),
    .O(net_42512_cascademuxed)
  );
  Span4Mux_v1 t5710 (
    .I(seg_25_13_sp4_h_l_45_84416),
    .O(seg_25_12_sp4_v_b_21_95683)
  );
  Span4Mux_h4 t5711 (
    .I(seg_21_13_sp4_h_l_45_69723),
    .O(seg_25_13_sp4_h_l_45_84416)
  );
  Span4Mux_h4 t5712 (
    .I(seg_17_13_sp4_v_b_2_65528),
    .O(seg_21_13_sp4_h_l_45_69723)
  );
  LocalMux t5713 (
    .I(seg_25_11_sp4_v_b_30_95681),
    .O(seg_25_11_local_g2_6_100172)
  );
  Span4Mux_v2 t5714 (
    .I(seg_25_13_sp4_h_l_43_84414),
    .O(seg_25_11_sp4_v_b_30_95681)
  );
  Span4Mux_h4 t5715 (
    .I(seg_21_13_sp4_h_l_47_69715),
    .O(seg_25_13_sp4_h_l_43_84414)
  );
  Span4Mux_h4 t5716 (
    .I(seg_17_13_sp4_v_b_4_65530),
    .O(seg_21_13_sp4_h_l_47_69715)
  );
  LocalMux t5717 (
    .I(seg_25_12_sp4_v_b_19_95681),
    .O(seg_25_12_local_g1_3_100311)
  );
  Span4Mux_v1 t5718 (
    .I(seg_25_13_sp4_h_l_43_84414),
    .O(seg_25_12_sp4_v_b_19_95681)
  );
  LocalMux t5719 (
    .I(seg_25_11_sp4_v_b_27_95676),
    .O(seg_25_11_local_g2_3_100169)
  );
  CascadeMux t572 (
    .I(net_42617),
    .O(net_42617_cascademuxed)
  );
  Span4Mux_v2 t5720 (
    .I(seg_25_13_sp4_h_l_38_84411),
    .O(seg_25_11_sp4_v_b_27_95676)
  );
  Span4Mux_h4 t5721 (
    .I(seg_21_13_sp4_h_l_37_69713),
    .O(seg_25_13_sp4_h_l_38_84411)
  );
  Span4Mux_h4 t5722 (
    .I(seg_17_13_sp4_v_b_6_65532),
    .O(seg_21_13_sp4_h_l_37_69713)
  );
  LocalMux t5723 (
    .I(seg_25_12_sp4_v_b_14_95676),
    .O(seg_25_12_local_g1_6_100314)
  );
  Span4Mux_v1 t5724 (
    .I(seg_25_13_sp4_h_l_38_84411),
    .O(seg_25_12_sp4_v_b_14_95676)
  );
  LocalMux t5725 (
    .I(seg_17_12_neigh_op_bnl_1_61671),
    .O(seg_17_12_local_g3_1_69521)
  );
  LocalMux t5726 (
    .I(seg_17_12_neigh_op_bnl_3_61673),
    .O(seg_17_12_local_g2_3_69515)
  );
  LocalMux t5727 (
    .I(seg_17_11_neigh_op_lft_5_61675),
    .O(seg_17_11_local_g0_5_69378)
  );
  LocalMux t5728 (
    .I(seg_15_11_neigh_op_rgt_6_61676),
    .O(seg_15_11_local_g2_6_61733)
  );
  LocalMux t5729 (
    .I(seg_15_11_neigh_op_rgt_7_61677),
    .O(seg_15_11_local_g2_7_61734)
  );
  CascadeMux t573 (
    .I(net_42635),
    .O(net_42635_cascademuxed)
  );
  LocalMux t5730 (
    .I(seg_16_31_span12_vert_2_66741),
    .O(seg_16_31_local_g1_2_68025)
  );
  Span12Mux_v11 t5731 (
    .I(seg_16_20_sp12_v_b_1_65265),
    .O(seg_16_31_span12_vert_2_66741)
  );
  LocalMux t5732 (
    .I(seg_16_31_span12_vert_6_66987),
    .O(seg_16_31_local_g0_6_68021)
  );
  Span12Mux_v9 t5733 (
    .I(seg_16_22_sp12_v_b_1_65511),
    .O(seg_16_31_span12_vert_6_66987)
  );
  LocalMux t5734 (
    .I(seg_18_0_span4_vert_24_68230),
    .O(seg_18_0_local_g1_0_71884)
  );
  Span4Mux_v3 t5735 (
    .I(seg_18_3_sp4_v_t_44_68626),
    .O(seg_18_0_span4_vert_24_68230)
  );
  Span4Mux_v4 t5736 (
    .I(seg_18_7_sp4_v_t_43_69117),
    .O(seg_18_3_sp4_v_t_44_68626)
  );
  Span4Mux_v4 t5737 (
    .I(seg_18_11_sp4_h_l_37_57975),
    .O(seg_18_7_sp4_v_t_43_69117)
  );
  LocalMux t5738 (
    .I(seg_18_31_span4_horz_r_5_71863),
    .O(seg_18_31_local_g0_5_75682)
  );
  IoSpan4Mux t5739 (
    .I(seg_17_31_span4_vert_7_67745),
    .O(seg_18_31_span4_horz_r_5_71863)
  );
  CascadeMux t574 (
    .I(net_42851),
    .O(net_42851_cascademuxed)
  );
  Span4Mux_v4 t5740 (
    .I(seg_17_27_sp4_v_b_7_67253),
    .O(seg_17_31_span4_vert_7_67745)
  );
  Span4Mux_v4 t5741 (
    .I(seg_17_23_sp4_v_b_4_66760),
    .O(seg_17_27_sp4_v_b_7_67253)
  );
  Span4Mux_v4 t5742 (
    .I(seg_17_19_sp4_v_b_1_66263),
    .O(seg_17_23_sp4_v_b_4_66760)
  );
  Span4Mux_v4 t5743 (
    .I(seg_17_15_sp4_v_b_1_65771),
    .O(seg_17_19_sp4_v_b_1_66263)
  );
  Span4Mux_v4 t5744 (
    .I(seg_17_11_sp4_h_l_36_54146),
    .O(seg_17_15_sp4_v_b_1_65771)
  );
  LocalMux t5745 (
    .I(seg_18_11_sp4_h_r_32_65646),
    .O(seg_18_11_local_g2_0_73220)
  );
  LocalMux t5746 (
    .I(seg_18_12_sp4_h_r_15_69594),
    .O(seg_18_12_local_g1_7_73342)
  );
  Span4Mux_h1 t5747 (
    .I(seg_17_12_sp4_v_b_8_65411),
    .O(seg_18_12_sp4_h_r_15_69594)
  );
  LocalMux t5748 (
    .I(seg_8_0_span4_vert_36_29935),
    .O(seg_8_0_local_g0_4_33572)
  );
  Span4Mux_v4 t5749 (
    .I(seg_8_4_sp4_h_r_1_34130),
    .O(seg_8_0_span4_vert_36_29935)
  );
  CascadeMux t575 (
    .I(net_42980),
    .O(net_42980_cascademuxed)
  );
  Span4Mux_h4 t5750 (
    .I(seg_12_4_sp4_h_r_10_49455),
    .O(seg_8_4_sp4_h_r_1_34130)
  );
  Span4Mux_h4 t5751 (
    .I(seg_16_4_sp4_v_t_41_61084),
    .O(seg_12_4_sp4_h_r_10_49455)
  );
  Span4Mux_v4 t5752 (
    .I(seg_16_8_sp4_v_t_36_61571),
    .O(seg_16_4_sp4_v_t_41_61084)
  );
  LocalMux t5753 (
    .I(seg_16_0_span4_vert_43_60589),
    .O(seg_16_0_local_g1_3_64225)
  );
  Span4Mux_v4 t5754 (
    .I(seg_16_4_sp4_v_t_43_61086),
    .O(seg_16_0_span4_vert_43_60589)
  );
  Span4Mux_v4 t5755 (
    .I(seg_16_8_sp4_v_t_38_61573),
    .O(seg_16_4_sp4_v_t_43_61086)
  );
  LocalMux t5756 (
    .I(seg_20_12_sp4_h_r_20_77010),
    .O(seg_20_12_local_g0_4_80362)
  );
  Span4Mux_h1 t5757 (
    .I(seg_19_12_sp4_h_l_36_61929),
    .O(seg_20_12_sp4_h_r_20_77010)
  );
  LocalMux t5758 (
    .I(seg_14_18_sp4_r_v_b_35_58735),
    .O(seg_14_18_local_g2_3_58761)
  );
  Span4Mux_v2 t5759 (
    .I(seg_15_16_sp4_v_b_3_58235),
    .O(seg_14_18_sp4_r_v_b_35_58735)
  );
  CascadeMux t576 (
    .I(net_43085),
    .O(net_43085_cascademuxed)
  );
  Span4Mux_v4 t5760 (
    .I(seg_15_12_sp4_h_r_9_61939),
    .O(seg_15_16_sp4_v_b_3_58235)
  );
  LocalMux t5761 (
    .I(seg_11_12_sp4_h_r_15_42779),
    .O(seg_11_12_local_g0_7_46519)
  );
  Span4Mux_h3 t5762 (
    .I(seg_14_12_sp4_h_r_6_58106),
    .O(seg_11_12_sp4_h_r_15_42779)
  );
  LocalMux t5763 (
    .I(seg_13_8_sp4_h_r_19_49953),
    .O(seg_13_8_local_g0_3_53685)
  );
  Span4Mux_h3 t5764 (
    .I(seg_16_8_sp4_v_t_43_61578),
    .O(seg_13_8_sp4_h_r_19_49953)
  );
  LocalMux t5765 (
    .I(seg_15_13_neigh_op_rgt_1_61917),
    .O(seg_15_13_local_g3_1_61982)
  );
  LocalMux t5766 (
    .I(seg_15_13_neigh_op_rgt_2_61918),
    .O(seg_15_13_local_g2_2_61975)
  );
  LocalMux t5767 (
    .I(seg_15_13_neigh_op_rgt_3_61919),
    .O(seg_15_13_local_g2_3_61976)
  );
  LocalMux t5768 (
    .I(seg_15_13_neigh_op_rgt_4_61920),
    .O(seg_15_13_local_g3_4_61985)
  );
  LocalMux t5769 (
    .I(seg_15_13_neigh_op_rgt_5_61921),
    .O(seg_15_13_local_g3_5_61986)
  );
  CascadeMux t577 (
    .I(net_43097),
    .O(net_43097_cascademuxed)
  );
  LocalMux t5770 (
    .I(seg_15_13_neigh_op_rgt_6_61922),
    .O(seg_15_13_local_g3_6_61987)
  );
  LocalMux t5771 (
    .I(seg_13_14_sp4_h_r_7_54523),
    .O(seg_13_14_local_g0_7_54427)
  );
  Span4Mux_h4 t5772 (
    .I(seg_17_14_sp4_v_b_2_65651),
    .O(seg_13_14_sp4_h_r_7_54523)
  );
  LocalMux t5773 (
    .I(seg_15_11_sp4_h_r_31_54154),
    .O(seg_15_11_local_g3_7_61742)
  );
  Span4Mux_h2 t5774 (
    .I(seg_17_11_sp4_v_t_42_65777),
    .O(seg_15_11_sp4_h_r_31_54154)
  );
  LocalMux t5775 (
    .I(seg_16_18_sp4_r_v_b_14_66265),
    .O(seg_16_18_local_g2_6_66425)
  );
  Span4Mux_v3 t5776 (
    .I(seg_17_15_sp4_v_b_7_65777),
    .O(seg_16_18_sp4_r_v_b_14_66265)
  );
  LocalMux t5777 (
    .I(seg_17_13_neigh_op_tnl_1_62040),
    .O(seg_17_13_local_g3_1_69644)
  );
  LocalMux t5778 (
    .I(seg_17_13_neigh_op_tnl_2_62041),
    .O(seg_17_13_local_g2_2_69637)
  );
  LocalMux t5779 (
    .I(seg_17_13_neigh_op_tnl_3_62042),
    .O(seg_17_13_local_g3_3_69646)
  );
  CascadeMux t578 (
    .I(net_43109),
    .O(net_43109_cascademuxed)
  );
  LocalMux t5780 (
    .I(seg_17_13_neigh_op_tnl_4_62043),
    .O(seg_17_13_local_g2_4_69639)
  );
  LocalMux t5781 (
    .I(seg_17_13_neigh_op_tnl_5_62044),
    .O(seg_17_13_local_g3_5_69648)
  );
  LocalMux t5782 (
    .I(seg_17_13_neigh_op_tnl_6_62045),
    .O(seg_17_13_local_g2_6_69641)
  );
  LocalMux t5783 (
    .I(seg_17_13_neigh_op_tnl_7_62046),
    .O(seg_17_13_local_g3_7_69650)
  );
  LocalMux t5784 (
    .I(seg_17_14_neigh_op_tnl_0_62162),
    .O(seg_17_14_local_g2_0_69758)
  );
  LocalMux t5785 (
    .I(seg_16_14_neigh_op_top_1_62163),
    .O(seg_16_14_local_g0_1_65912)
  );
  LocalMux t5786 (
    .I(seg_16_14_neigh_op_top_2_62164),
    .O(seg_16_14_local_g0_2_65913)
  );
  LocalMux t5787 (
    .I(seg_16_15_lutff_4_out_62166),
    .O(seg_16_15_local_g2_4_66054)
  );
  LocalMux t5788 (
    .I(seg_15_14_neigh_op_tnr_5_62167),
    .O(seg_15_14_local_g3_5_62109)
  );
  LocalMux t5789 (
    .I(seg_15_15_neigh_op_rgt_6_62168),
    .O(seg_15_15_local_g3_6_62233)
  );
  CascadeMux t579 (
    .I(net_43226),
    .O(net_43226_cascademuxed)
  );
  LocalMux t5790 (
    .I(seg_16_14_neigh_op_top_7_62169),
    .O(seg_16_14_local_g1_7_65926)
  );
  LocalMux t5791 (
    .I(seg_18_15_sp4_h_r_34_66130),
    .O(seg_18_15_local_g3_2_73722)
  );
  LocalMux t5792 (
    .I(seg_18_15_sp4_h_r_36_62298),
    .O(seg_18_15_local_g3_4_73724)
  );
  LocalMux t5793 (
    .I(seg_18_16_sp4_v_b_37_70095),
    .O(seg_18_16_local_g3_5_73848)
  );
  Span4Mux_v1 t5794 (
    .I(seg_18_15_sp4_h_l_37_58467),
    .O(seg_18_16_sp4_v_b_37_70095)
  );
  LocalMux t5795 (
    .I(seg_17_12_sp4_v_b_46_65781),
    .O(seg_17_12_local_g3_6_69526)
  );
  LocalMux t5796 (
    .I(seg_16_13_sp4_v_b_46_62073),
    .O(seg_16_13_local_g2_6_65810)
  );
  LocalMux t5797 (
    .I(seg_15_16_neigh_op_rgt_0_62285),
    .O(seg_15_16_local_g2_0_62342)
  );
  LocalMux t5798 (
    .I(seg_15_16_neigh_op_rgt_1_62286),
    .O(seg_15_16_local_g3_1_62351)
  );
  LocalMux t5799 (
    .I(seg_17_15_neigh_op_tnl_2_62287),
    .O(seg_17_15_local_g3_2_69891)
  );
  CascadeMux t58 (
    .I(net_11324),
    .O(net_11324_cascademuxed)
  );
  CascadeMux t580 (
    .I(net_43331),
    .O(net_43331_cascademuxed)
  );
  LocalMux t5800 (
    .I(seg_16_16_lutff_3_out_62288),
    .O(seg_16_16_local_g2_3_66176)
  );
  LocalMux t5801 (
    .I(seg_17_15_neigh_op_tnl_3_62288),
    .O(seg_17_15_local_g3_3_69892)
  );
  LocalMux t5802 (
    .I(seg_16_16_lutff_4_out_62289),
    .O(seg_16_16_local_g0_4_66161)
  );
  LocalMux t5803 (
    .I(seg_15_16_neigh_op_rgt_6_62291),
    .O(seg_15_16_local_g3_6_62356)
  );
  LocalMux t5804 (
    .I(seg_16_15_neigh_op_top_7_62292),
    .O(seg_16_15_local_g1_7_66049)
  );
  LocalMux t5805 (
    .I(seg_16_16_lutff_7_out_62292),
    .O(seg_16_16_local_g2_7_66180)
  );
  LocalMux t5806 (
    .I(seg_14_16_sp4_h_r_8_58600),
    .O(seg_14_16_local_g0_0_58496)
  );
  LocalMux t5807 (
    .I(seg_14_16_sp4_h_r_10_58592),
    .O(seg_14_16_local_g1_2_58506)
  );
  LocalMux t5808 (
    .I(seg_14_16_sp4_h_r_20_54771),
    .O(seg_14_16_local_g0_4_58500)
  );
  LocalMux t5809 (
    .I(seg_18_16_sp4_h_r_32_66261),
    .O(seg_18_16_local_g2_0_73835)
  );
  CascadeMux t581 (
    .I(net_43343),
    .O(net_43343_cascademuxed)
  );
  LocalMux t5810 (
    .I(seg_18_16_sp4_h_r_16_70089),
    .O(seg_18_16_local_g0_0_73819)
  );
  Span4Mux_h1 t5811 (
    .I(seg_17_16_sp4_v_b_11_65904),
    .O(seg_18_16_sp4_h_r_16_70089)
  );
  LocalMux t5812 (
    .I(seg_16_16_neigh_op_top_0_62408),
    .O(seg_16_16_local_g1_0_66165)
  );
  LocalMux t5813 (
    .I(seg_16_17_lutff_1_out_62409),
    .O(seg_16_17_local_g3_1_66305)
  );
  LocalMux t5814 (
    .I(seg_15_16_neigh_op_tnr_2_62410),
    .O(seg_15_16_local_g3_2_62352)
  );
  LocalMux t5815 (
    .I(seg_15_17_neigh_op_rgt_3_62411),
    .O(seg_15_17_local_g2_3_62468)
  );
  LocalMux t5816 (
    .I(seg_16_17_lutff_3_out_62411),
    .O(seg_16_17_local_g2_3_66299)
  );
  LocalMux t5817 (
    .I(seg_16_17_lutff_4_out_62412),
    .O(seg_16_17_local_g3_4_66308)
  );
  LocalMux t5818 (
    .I(seg_16_17_lutff_5_out_62413),
    .O(seg_16_17_local_g1_5_66293)
  );
  LocalMux t5819 (
    .I(seg_16_17_lutff_6_out_62414),
    .O(seg_16_17_local_g3_6_66310)
  );
  CascadeMux t582 (
    .I(net_43367),
    .O(net_43367_cascademuxed)
  );
  LocalMux t5820 (
    .I(seg_18_16_sp4_r_v_b_14_73681),
    .O(seg_18_16_local_g2_6_73841)
  );
  Span4Mux_v1 t5821 (
    .I(seg_19_17_sp4_h_l_38_62548),
    .O(seg_18_16_sp4_r_v_b_14_73681)
  );
  LocalMux t5822 (
    .I(seg_14_17_sp4_h_r_14_54888),
    .O(seg_14_17_local_g1_6_58633)
  );
  LocalMux t5823 (
    .I(seg_17_15_sp4_v_b_37_66141),
    .O(seg_17_15_local_g3_5_69894)
  );
  LocalMux t5824 (
    .I(seg_17_15_sp4_v_b_27_66019),
    .O(seg_17_15_local_g2_3_69884)
  );
  LocalMux t5825 (
    .I(seg_18_16_sp4_h_r_19_70090),
    .O(seg_18_16_local_g1_3_73830)
  );
  Span4Mux_h1 t5826 (
    .I(seg_17_16_sp4_v_t_43_66393),
    .O(seg_18_16_sp4_h_r_19_70090)
  );
  LocalMux t5827 (
    .I(seg_17_15_sp4_v_b_33_66025),
    .O(seg_17_15_local_g2_1_69882)
  );
  LocalMux t5828 (
    .I(seg_16_15_sp4_v_b_24_62187),
    .O(seg_16_15_local_g2_0_66050)
  );
  LocalMux t5829 (
    .I(seg_14_16_sp4_h_r_31_50938),
    .O(seg_14_16_local_g3_7_58527)
  );
  CascadeMux t583 (
    .I(net_43454),
    .O(net_43454_cascademuxed)
  );
  Span4Mux_h2 t5830 (
    .I(seg_16_16_sp4_v_t_36_62555),
    .O(seg_14_16_sp4_h_r_31_50938)
  );
  LocalMux t5831 (
    .I(seg_14_13_sp4_h_r_24_50560),
    .O(seg_14_13_local_g2_0_58143)
  );
  Span4Mux_h2 t5832 (
    .I(seg_16_13_sp4_v_t_43_62193),
    .O(seg_14_13_sp4_h_r_24_50560)
  );
  LocalMux t5833 (
    .I(seg_16_13_sp12_v_b_11_65020),
    .O(seg_16_13_local_g3_3_65815)
  );
  LocalMux t5834 (
    .I(seg_3_1_sp4_h_r_13_11369),
    .O(seg_3_1_local_g1_5_15115)
  );
  Span4Mux_h3 t5835 (
    .I(seg_6_1_sp4_h_r_9_26682),
    .O(seg_3_1_sp4_h_r_13_11369)
  );
  Span4Mux_h4 t5836 (
    .I(seg_10_1_sp4_h_r_1_41387),
    .O(seg_6_1_sp4_h_r_9_26682)
  );
  Span4Mux_h4 t5837 (
    .I(seg_14_1_sp4_v_b_1_52892),
    .O(seg_10_1_sp4_h_r_1_41387)
  );
  IoSpan4Mux t5838 (
    .I(seg_14_0_span4_horz_r_0_56601),
    .O(seg_14_1_sp4_v_b_1_52892)
  );
  LocalMux t5839 (
    .I(seg_4_2_sp4_r_v_b_13_19060),
    .O(seg_4_2_local_g2_5_19117)
  );
  CascadeMux t584 (
    .I(net_43460),
    .O(net_43460_cascademuxed)
  );
  Span4Mux_v1 t5840 (
    .I(seg_5_3_sp4_h_r_0_23144),
    .O(seg_4_2_sp4_r_v_b_13_19060)
  );
  Span4Mux_h4 t5841 (
    .I(seg_9_3_sp4_h_r_4_37843),
    .O(seg_5_3_sp4_h_r_0_23144)
  );
  Span4Mux_h4 t5842 (
    .I(seg_13_3_sp4_h_r_8_53171),
    .O(seg_9_3_sp4_h_r_4_37843)
  );
  Span4Mux_h4 t5843 (
    .I(seg_17_3_sp4_v_b_8_64408),
    .O(seg_13_3_sp4_h_r_8_53171)
  );
  LocalMux t5844 (
    .I(seg_20_6_sp4_r_v_b_5_79361),
    .O(seg_20_6_local_g1_5_79633)
  );
  Span4Mux_v4 t5845 (
    .I(seg_21_2_sp4_h_l_37_68360),
    .O(seg_20_6_sp4_r_v_b_5_79361)
  );
  LocalMux t5846 (
    .I(seg_20_6_sp4_v_b_3_76095),
    .O(seg_20_6_local_g1_3_79631)
  );
  Span4Mux_v4 t5847 (
    .I(seg_20_2_sp4_h_l_38_64534),
    .O(seg_20_6_sp4_v_b_3_76095)
  );
  LocalMux t5848 (
    .I(seg_17_3_lutff_0_out_64517),
    .O(seg_17_3_local_g3_0_68413)
  );
  LocalMux t5849 (
    .I(seg_18_4_neigh_op_bnl_1_64518),
    .O(seg_18_4_local_g2_1_72360)
  );
  CascadeMux t585 (
    .I(net_43466),
    .O(net_43466_cascademuxed)
  );
  LocalMux t5850 (
    .I(seg_16_4_neigh_op_bnr_3_64520),
    .O(seg_16_4_local_g1_3_64692)
  );
  LocalMux t5851 (
    .I(seg_16_4_neigh_op_bnr_4_64521),
    .O(seg_16_4_local_g1_4_64693)
  );
  LocalMux t5852 (
    .I(seg_15_3_sp4_h_r_12_56992),
    .O(seg_15_3_local_g0_4_60731)
  );
  LocalMux t5853 (
    .I(seg_16_4_neigh_op_rgt_0_64640),
    .O(seg_16_4_local_g3_0_64705)
  );
  LocalMux t5854 (
    .I(seg_16_4_neigh_op_rgt_1_64641),
    .O(seg_16_4_local_g2_1_64698)
  );
  LocalMux t5855 (
    .I(seg_16_4_neigh_op_rgt_3_64643),
    .O(seg_16_4_local_g2_3_64700)
  );
  LocalMux t5856 (
    .I(seg_16_4_neigh_op_rgt_4_64644),
    .O(seg_16_4_local_g2_4_64701)
  );
  LocalMux t5857 (
    .I(seg_16_4_neigh_op_rgt_5_64645),
    .O(seg_16_4_local_g2_5_64702)
  );
  LocalMux t5858 (
    .I(seg_16_4_neigh_op_rgt_6_64646),
    .O(seg_16_4_local_g2_6_64703)
  );
  LocalMux t5859 (
    .I(seg_16_4_neigh_op_rgt_7_64647),
    .O(seg_16_4_local_g3_7_64712)
  );
  CascadeMux t586 (
    .I(net_43478),
    .O(net_43478_cascademuxed)
  );
  LocalMux t5860 (
    .I(seg_18_4_sp4_v_b_5_68248),
    .O(seg_18_4_local_g1_5_72356)
  );
  LocalMux t5861 (
    .I(seg_16_4_neigh_op_tnr_0_64763),
    .O(seg_16_4_local_g2_0_64697)
  );
  LocalMux t5862 (
    .I(seg_16_5_neigh_op_rgt_0_64763),
    .O(seg_16_5_local_g2_0_64820)
  );
  LocalMux t5863 (
    .I(seg_16_5_neigh_op_rgt_1_64764),
    .O(seg_16_5_local_g3_1_64829)
  );
  LocalMux t5864 (
    .I(seg_16_5_neigh_op_rgt_2_64765),
    .O(seg_16_5_local_g2_2_64822)
  );
  LocalMux t5865 (
    .I(seg_16_5_neigh_op_rgt_3_64766),
    .O(seg_16_5_local_g2_3_64823)
  );
  LocalMux t5866 (
    .I(seg_18_4_neigh_op_tnl_5_64768),
    .O(seg_18_4_local_g2_5_72364)
  );
  LocalMux t5867 (
    .I(seg_18_6_neigh_op_bnl_5_64768),
    .O(seg_18_6_local_g3_5_72618)
  );
  LocalMux t5868 (
    .I(seg_16_4_neigh_op_tnr_6_64769),
    .O(seg_16_4_local_g3_6_64711)
  );
  LocalMux t5869 (
    .I(seg_16_5_neigh_op_rgt_6_64769),
    .O(seg_16_5_local_g2_6_64826)
  );
  CascadeMux t587 (
    .I(net_43484),
    .O(net_43484_cascademuxed)
  );
  LocalMux t5870 (
    .I(seg_16_5_neigh_op_rgt_7_64770),
    .O(seg_16_5_local_g3_7_64835)
  );
  LocalMux t5871 (
    .I(seg_16_5_neigh_op_tnr_2_64888),
    .O(seg_16_5_local_g3_2_64830)
  );
  LocalMux t5872 (
    .I(seg_16_7_neigh_op_bnr_4_64890),
    .O(seg_16_7_local_g0_4_65054)
  );
  LocalMux t5873 (
    .I(seg_17_6_lutff_5_out_64891),
    .O(seg_17_6_local_g2_5_68779)
  );
  LocalMux t5874 (
    .I(seg_16_5_neigh_op_tnr_6_64892),
    .O(seg_16_5_local_g3_6_64834)
  );
  LocalMux t5875 (
    .I(seg_12_6_sp4_h_r_11_49702),
    .O(seg_12_6_local_g1_3_49616)
  );
  Span4Mux_h4 t5876 (
    .I(seg_16_6_sp4_h_r_3_65026),
    .O(seg_12_6_sp4_h_r_11_49702)
  );
  LocalMux t5877 (
    .I(seg_17_7_lutff_7_out_65016),
    .O(seg_17_7_local_g0_7_68888)
  );
  LocalMux t5878 (
    .I(seg_14_3_sp4_h_r_11_56994),
    .O(seg_14_3_local_g0_3_56900)
  );
  Span4Mux_h0 t5879 (
    .I(seg_14_3_sp4_v_t_46_53306),
    .O(seg_14_3_sp4_h_r_11_56994)
  );
  CascadeMux t588 (
    .I(net_43496),
    .O(net_43496_cascademuxed)
  );
  Span4Mux_v4 t5880 (
    .I(seg_14_7_sp4_h_r_11_57486),
    .O(seg_14_3_sp4_v_t_46_53306)
  );
  LocalMux t5881 (
    .I(seg_12_1_sp4_r_v_b_45_49100),
    .O(seg_12_1_local_g3_5_48979)
  );
  Span4Mux_v3 t5882 (
    .I(seg_13_4_sp4_h_r_3_53289),
    .O(seg_12_1_sp4_r_v_b_45_49100)
  );
  Span4Mux_h4 t5883 (
    .I(seg_17_4_sp4_v_t_38_64912),
    .O(seg_13_4_sp4_h_r_3_53289)
  );
  LocalMux t5884 (
    .I(seg_13_3_sp4_v_b_21_49100),
    .O(seg_13_3_local_g1_5_53080)
  );
  Span4Mux_v1 t5885 (
    .I(seg_13_4_sp4_h_r_3_53289),
    .O(seg_13_3_sp4_v_b_21_49100)
  );
  LocalMux t5886 (
    .I(seg_13_4_sp4_h_r_3_53289),
    .O(seg_13_4_local_g0_3_53193)
  );
  LocalMux t5887 (
    .I(seg_13_8_sp4_h_r_30_46122),
    .O(seg_13_8_local_g3_6_53712)
  );
  Span4Mux_h2 t5888 (
    .I(seg_15_8_sp4_h_r_10_61438),
    .O(seg_13_8_sp4_h_r_30_46122)
  );
  LocalMux t5889 (
    .I(seg_13_8_sp4_r_v_b_1_53419),
    .O(seg_13_8_local_g1_1_53691)
  );
  CascadeMux t589 (
    .I(net_43583),
    .O(net_43583_cascademuxed)
  );
  Span4Mux_v1 t5890 (
    .I(seg_14_8_sp4_h_r_1_57607),
    .O(seg_13_8_sp4_r_v_b_1_53419)
  );
  LocalMux t5891 (
    .I(seg_13_8_sp4_r_v_b_9_53427),
    .O(seg_13_8_local_g2_1_53699)
  );
  Span4Mux_v1 t5892 (
    .I(seg_14_8_sp4_h_r_9_57617),
    .O(seg_13_8_sp4_r_v_b_9_53427)
  );
  LocalMux t5893 (
    .I(seg_16_9_neigh_op_rgt_7_65262),
    .O(seg_16_9_local_g3_7_65327)
  );
  LocalMux t5894 (
    .I(seg_17_4_sp4_v_b_22_64551),
    .O(seg_17_4_local_g1_6_68526)
  );
  Span4Mux_v1 t5895 (
    .I(seg_17_5_sp4_v_t_45_65042),
    .O(seg_17_4_sp4_v_b_22_64551)
  );
  LocalMux t5896 (
    .I(seg_17_11_neigh_op_bot_0_65378),
    .O(seg_17_11_local_g0_0_69373)
  );
  LocalMux t5897 (
    .I(seg_16_10_neigh_op_rgt_1_65379),
    .O(seg_16_10_local_g2_1_65436)
  );
  LocalMux t5898 (
    .I(seg_17_11_neigh_op_bot_1_65379),
    .O(seg_17_11_local_g0_1_69374)
  );
  LocalMux t5899 (
    .I(seg_18_9_neigh_op_tnl_2_65380),
    .O(seg_18_9_local_g2_2_72976)
  );
  CascadeMux t59 (
    .I(net_11336),
    .O(net_11336_cascademuxed)
  );
  CascadeMux t590 (
    .I(net_43619),
    .O(net_43619_cascademuxed)
  );
  LocalMux t5900 (
    .I(seg_18_10_neigh_op_lft_2_65380),
    .O(seg_18_10_local_g1_2_73091)
  );
  LocalMux t5901 (
    .I(seg_16_11_neigh_op_bnr_5_65383),
    .O(seg_16_11_local_g0_5_65547)
  );
  LocalMux t5902 (
    .I(seg_16_11_neigh_op_bnr_5_65383),
    .O(seg_16_11_local_g1_5_65555)
  );
  LocalMux t5903 (
    .I(seg_17_11_neigh_op_bot_5_65383),
    .O(seg_17_11_local_g1_5_69386)
  );
  LocalMux t5904 (
    .I(seg_17_10_lutff_7_out_65385),
    .O(seg_17_10_local_g1_7_69265)
  );
  LocalMux t5905 (
    .I(seg_10_10_sp12_h_r_1_42526),
    .O(seg_10_10_local_g1_1_42444)
  );
  LocalMux t5906 (
    .I(seg_15_12_sp4_v_b_30_57994),
    .O(seg_15_12_local_g3_6_61864)
  );
  Span4Mux_v2 t5907 (
    .I(seg_15_10_sp4_h_r_0_61682),
    .O(seg_15_12_sp4_v_b_30_57994)
  );
  LocalMux t5908 (
    .I(seg_15_13_sp4_v_b_19_57994),
    .O(seg_15_13_local_g1_3_61968)
  );
  Span4Mux_v3 t5909 (
    .I(seg_15_10_sp4_h_r_0_61682),
    .O(seg_15_13_sp4_v_b_19_57994)
  );
  LocalMux t5910 (
    .I(seg_11_5_sp4_v_b_19_41687),
    .O(seg_11_5_local_g0_3_45654)
  );
  Span4Mux_v1 t5911 (
    .I(seg_11_6_sp4_h_r_1_45869),
    .O(seg_11_5_sp4_v_b_19_41687)
  );
  Span4Mux_h4 t5912 (
    .I(seg_15_6_sp4_v_t_42_57501),
    .O(seg_11_6_sp4_h_r_1_45869)
  );
  Span4Mux_v4 t5913 (
    .I(seg_15_10_sp4_h_r_2_61686),
    .O(seg_15_6_sp4_v_t_42_57501)
  );
  LocalMux t5914 (
    .I(seg_18_7_sp4_v_b_46_68997),
    .O(seg_18_7_local_g3_6_72742)
  );
  LocalMux t5915 (
    .I(seg_18_8_sp4_v_b_35_68997),
    .O(seg_18_8_local_g2_3_72854)
  );
  LocalMux t5916 (
    .I(seg_7_6_sp4_h_r_27_23518),
    .O(seg_7_6_local_g3_3_30477)
  );
  Span4Mux_h2 t5917 (
    .I(seg_9_6_sp4_h_r_0_38206),
    .O(seg_7_6_sp4_h_r_27_23518)
  );
  Span4Mux_h4 t5918 (
    .I(seg_13_6_sp4_h_r_4_53536),
    .O(seg_9_6_sp4_h_r_0_38206)
  );
  Span4Mux_h4 t5919 (
    .I(seg_17_6_sp4_v_t_47_65167),
    .O(seg_13_6_sp4_h_r_4_53536)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t592 (
    .carryinitin(),
    .carryinitout(t591)
  );
  LocalMux t5920 (
    .I(seg_11_4_sp4_h_r_26_37964),
    .O(seg_11_4_local_g2_2_45546)
  );
  Span4Mux_h2 t5921 (
    .I(seg_13_4_sp4_h_r_11_53287),
    .O(seg_11_4_sp4_h_r_26_37964)
  );
  Span4Mux_h4 t5922 (
    .I(seg_17_4_sp4_v_t_40_64914),
    .O(seg_13_4_sp4_h_r_11_53287)
  );
  Span4Mux_v4 t5923 (
    .I(seg_17_8_sp4_v_t_39_65405),
    .O(seg_17_4_sp4_v_t_40_64914)
  );
  LocalMux t5924 (
    .I(seg_11_4_sp4_h_r_26_37964),
    .O(seg_11_4_local_g3_2_45554)
  );
  LocalMux t5925 (
    .I(seg_16_11_neigh_op_rgt_1_65502),
    .O(seg_16_11_local_g3_1_65567)
  );
  LocalMux t5926 (
    .I(seg_16_11_neigh_op_rgt_2_65503),
    .O(seg_16_11_local_g3_2_65568)
  );
  LocalMux t5927 (
    .I(seg_16_11_neigh_op_rgt_3_65504),
    .O(seg_16_11_local_g3_3_65569)
  );
  LocalMux t5928 (
    .I(seg_16_11_neigh_op_rgt_4_65505),
    .O(seg_16_11_local_g2_4_65562)
  );
  LocalMux t5929 (
    .I(seg_17_11_lutff_5_out_65506),
    .O(seg_17_11_local_g3_5_69402)
  );
  LocalMux t5930 (
    .I(seg_18_11_neigh_op_lft_6_65507),
    .O(seg_18_11_local_g0_6_73210)
  );
  LocalMux t5931 (
    .I(seg_18_11_neigh_op_lft_7_65508),
    .O(seg_18_11_local_g0_7_73211)
  );
  LocalMux t5932 (
    .I(seg_17_31_span4_vert_1_67739),
    .O(seg_17_31_local_g1_1_71855)
  );
  Sp12to4 t5933 (
    .I(seg_17_30_sp12_v_b_1_70326),
    .O(seg_17_31_span4_vert_1_67739)
  );
  Span12Mux_v12 t5934 (
    .I(seg_17_18_sp12_v_b_1_68850),
    .O(seg_17_30_sp12_v_b_1_70326)
  );
  LocalMux t5935 (
    .I(seg_21_0_span4_vert_36_79105),
    .O(seg_21_0_local_g1_4_82750)
  );
  Span4Mux_v4 t5936 (
    .I(seg_21_4_sp4_h_l_36_68607),
    .O(seg_21_0_span4_vert_36_79105)
  );
  Span4Mux_h4 t5937 (
    .I(seg_17_4_sp4_v_t_36_64910),
    .O(seg_21_4_sp4_h_l_36_68607)
  );
  Span4Mux_v4 t5938 (
    .I(seg_17_8_sp4_v_t_36_65402),
    .O(seg_17_4_sp4_v_t_36_64910)
  );
  LocalMux t5939 (
    .I(seg_17_11_neigh_op_top_0_65624),
    .O(seg_17_11_local_g1_0_69381)
  );
  CascadeMux t594 (
    .I(net_45178),
    .O(net_45178_cascademuxed)
  );
  LocalMux t5940 (
    .I(seg_18_12_neigh_op_lft_1_65625),
    .O(seg_18_12_local_g1_1_73336)
  );
  LocalMux t5941 (
    .I(seg_17_12_lutff_2_out_65626),
    .O(seg_17_12_local_g3_2_69522)
  );
  LocalMux t5942 (
    .I(seg_17_12_lutff_3_out_65627),
    .O(seg_17_12_local_g0_3_69499)
  );
  LocalMux t5943 (
    .I(seg_17_11_neigh_op_top_4_65628),
    .O(seg_17_11_local_g1_4_69385)
  );
  LocalMux t5944 (
    .I(seg_17_12_lutff_5_out_65629),
    .O(seg_17_12_local_g3_5_69525)
  );
  LocalMux t5945 (
    .I(seg_17_12_lutff_6_out_65630),
    .O(seg_17_12_local_g2_6_69518)
  );
  LocalMux t5946 (
    .I(seg_17_11_neigh_op_top_7_65631),
    .O(seg_17_11_local_g1_7_69388)
  );
  LocalMux t5947 (
    .I(seg_17_14_neigh_op_bot_2_65749),
    .O(seg_17_14_local_g0_2_69744)
  );
  LocalMux t5948 (
    .I(seg_17_14_neigh_op_bot_3_65750),
    .O(seg_17_14_local_g1_3_69753)
  );
  LocalMux t5949 (
    .I(seg_17_14_neigh_op_bot_4_65751),
    .O(seg_17_14_local_g1_4_69754)
  );
  CascadeMux t595 (
    .I(net_45317),
    .O(net_45317_cascademuxed)
  );
  LocalMux t5950 (
    .I(seg_17_14_neigh_op_bot_5_65752),
    .O(seg_17_14_local_g1_5_69755)
  );
  LocalMux t5951 (
    .I(seg_17_14_neigh_op_bot_6_65753),
    .O(seg_17_14_local_g1_6_69756)
  );
  LocalMux t5952 (
    .I(seg_17_17_sp4_v_b_8_66026),
    .O(seg_17_17_local_g1_0_70119)
  );
  Span4Mux_v4 t5953 (
    .I(seg_17_13_sp4_h_r_2_69717),
    .O(seg_17_17_sp4_v_b_8_66026)
  );
  LocalMux t5954 (
    .I(seg_18_14_neigh_op_lft_1_65871),
    .O(seg_18_14_local_g1_1_73582)
  );
  LocalMux t5955 (
    .I(seg_18_14_neigh_op_lft_2_65872),
    .O(seg_18_14_local_g0_2_73575)
  );
  LocalMux t5956 (
    .I(seg_18_14_neigh_op_lft_3_65873),
    .O(seg_18_14_local_g0_3_73576)
  );
  LocalMux t5957 (
    .I(seg_17_13_neigh_op_top_4_65874),
    .O(seg_17_13_local_g0_4_69623)
  );
  LocalMux t5958 (
    .I(seg_16_14_neigh_op_rgt_5_65875),
    .O(seg_16_14_local_g3_5_65940)
  );
  LocalMux t5959 (
    .I(seg_17_14_lutff_5_out_65875),
    .O(seg_17_14_local_g2_5_69763)
  );
  CascadeMux t596 (
    .I(net_45323),
    .O(net_45323_cascademuxed)
  );
  LocalMux t5960 (
    .I(seg_18_14_neigh_op_lft_6_65876),
    .O(seg_18_14_local_g1_6_73587)
  );
  LocalMux t5961 (
    .I(seg_16_15_neigh_op_bnr_7_65877),
    .O(seg_16_15_local_g0_7_66041)
  );
  LocalMux t5962 (
    .I(seg_17_17_sp4_v_b_19_66147),
    .O(seg_17_17_local_g0_3_70114)
  );
  Span4Mux_v3 t5963 (
    .I(seg_17_14_sp4_h_r_0_69836),
    .O(seg_17_17_sp4_v_b_19_66147)
  );
  LocalMux t5964 (
    .I(seg_17_17_sp4_v_b_5_66021),
    .O(seg_17_17_local_g1_5_70124)
  );
  LocalMux t5965 (
    .I(seg_16_14_neigh_op_tnr_0_65993),
    .O(seg_16_14_local_g3_0_65935)
  );
  LocalMux t5966 (
    .I(seg_16_15_neigh_op_rgt_1_65994),
    .O(seg_16_15_local_g2_1_66051)
  );
  LocalMux t5967 (
    .I(seg_18_15_neigh_op_lft_1_65994),
    .O(seg_18_15_local_g0_1_73697)
  );
  LocalMux t5968 (
    .I(seg_16_14_neigh_op_tnr_2_65995),
    .O(seg_16_14_local_g3_2_65937)
  );
  LocalMux t5969 (
    .I(seg_16_14_neigh_op_tnr_3_65996),
    .O(seg_16_14_local_g2_3_65930)
  );
  CascadeMux t597 (
    .I(net_45329),
    .O(net_45329_cascademuxed)
  );
  LocalMux t5970 (
    .I(seg_17_14_neigh_op_top_4_65997),
    .O(seg_17_14_local_g0_4_69746)
  );
  LocalMux t5971 (
    .I(seg_18_15_neigh_op_lft_4_65997),
    .O(seg_18_15_local_g0_4_73700)
  );
  LocalMux t5972 (
    .I(seg_18_16_neigh_op_bnl_4_65997),
    .O(seg_18_16_local_g2_4_73839)
  );
  LocalMux t5973 (
    .I(seg_16_15_neigh_op_rgt_5_65998),
    .O(seg_16_15_local_g3_5_66063)
  );
  LocalMux t5974 (
    .I(seg_18_15_neigh_op_lft_5_65998),
    .O(seg_18_15_local_g0_5_73701)
  );
  LocalMux t5975 (
    .I(seg_16_15_neigh_op_rgt_6_65999),
    .O(seg_16_15_local_g3_6_66064)
  );
  LocalMux t5976 (
    .I(seg_18_15_neigh_op_lft_6_65999),
    .O(seg_18_15_local_g0_6_73702)
  );
  LocalMux t5977 (
    .I(seg_16_14_neigh_op_tnr_7_66000),
    .O(seg_16_14_local_g2_7_65934)
  );
  LocalMux t5978 (
    .I(seg_17_14_neigh_op_top_7_66000),
    .O(seg_17_14_local_g1_7_69757)
  );
  LocalMux t5979 (
    .I(seg_18_15_neigh_op_lft_7_66000),
    .O(seg_18_15_local_g0_7_73703)
  );
  CascadeMux t598 (
    .I(net_45347),
    .O(net_45347_cascademuxed)
  );
  LocalMux t5980 (
    .I(seg_18_16_neigh_op_bnl_7_66000),
    .O(seg_18_16_local_g3_7_73850)
  );
  LocalMux t5981 (
    .I(seg_18_15_sp4_h_r_17_69965),
    .O(seg_18_15_local_g1_1_73705)
  );
  LocalMux t5982 (
    .I(seg_18_13_sp4_v_b_27_69604),
    .O(seg_18_13_local_g3_3_73477)
  );
  LocalMux t5983 (
    .I(seg_18_13_sp4_v_b_33_69610),
    .O(seg_18_13_local_g3_1_73475)
  );
  LocalMux t5984 (
    .I(seg_17_10_sp4_v_b_28_65407),
    .O(seg_17_10_local_g2_4_69270)
  );
  Span4Mux_v2 t5985 (
    .I(seg_17_12_sp4_v_t_36_65894),
    .O(seg_17_10_sp4_v_b_28_65407)
  );
  LocalMux t5986 (
    .I(seg_17_17_neigh_op_bot_1_66117),
    .O(seg_17_17_local_g1_1_70120)
  );
  LocalMux t5987 (
    .I(seg_17_14_sp4_v_b_34_65905),
    .O(seg_17_14_local_g3_2_69768)
  );
  LocalMux t5988 (
    .I(seg_17_14_sp4_v_b_36_66017),
    .O(seg_17_14_local_g3_4_69770)
  );
  LocalMux t5989 (
    .I(seg_17_14_sp4_v_b_28_65899),
    .O(seg_17_14_local_g2_4_69762)
  );
  CascadeMux t599 (
    .I(net_45353),
    .O(net_45353_cascademuxed)
  );
  LocalMux t5990 (
    .I(seg_17_14_sp4_v_b_30_65901),
    .O(seg_17_14_local_g3_6_69772)
  );
  LocalMux t5991 (
    .I(seg_17_14_sp4_v_b_32_65903),
    .O(seg_17_14_local_g3_0_69766)
  );
  LocalMux t5992 (
    .I(seg_18_16_neigh_op_tnl_0_66239),
    .O(seg_18_16_local_g3_0_73843)
  );
  LocalMux t5993 (
    .I(seg_17_17_lutff_3_out_66242),
    .O(seg_17_17_local_g3_3_70138)
  );
  LocalMux t5994 (
    .I(seg_17_18_neigh_op_bot_4_66243),
    .O(seg_17_18_local_g0_4_70238)
  );
  LocalMux t5995 (
    .I(seg_17_17_lutff_5_out_66244),
    .O(seg_17_17_local_g0_5_70116)
  );
  LocalMux t5996 (
    .I(seg_15_16_sp4_r_v_b_14_62188),
    .O(seg_15_16_local_g2_6_62348)
  );
  Span4Mux_v1 t5997 (
    .I(seg_16_17_sp4_h_r_3_66379),
    .O(seg_15_16_sp4_r_v_b_14_62188)
  );
  LocalMux t5998 (
    .I(seg_15_16_sp4_v_b_16_58360),
    .O(seg_15_16_local_g0_0_62326)
  );
  Span4Mux_v1 t5999 (
    .I(seg_15_17_sp4_h_r_0_62543),
    .O(seg_15_16_sp4_v_b_16_58360)
  );
  CascadeMux t6 (
    .I(net_6792),
    .O(net_6792_cascademuxed)
  );
  CascadeMux t60 (
    .I(net_11348),
    .O(net_11348_cascademuxed)
  );
  CascadeMux t600 (
    .I(net_45440),
    .O(net_45440_cascademuxed)
  );
  LocalMux t6000 (
    .I(seg_15_17_sp4_h_r_16_58720),
    .O(seg_15_17_local_g0_0_62449)
  );
  LocalMux t6001 (
    .I(seg_14_17_sp4_h_r_11_58716),
    .O(seg_14_17_local_g1_3_58630)
  );
  LocalMux t6002 (
    .I(seg_18_14_sp4_h_r_0_73667),
    .O(seg_18_14_local_g0_0_73573)
  );
  Span4Mux_h0 t6003 (
    .I(seg_18_14_sp4_v_t_37_69972),
    .O(seg_18_14_sp4_h_r_0_73667)
  );
  LocalMux t6004 (
    .I(seg_17_15_sp4_r_v_b_27_69850),
    .O(seg_17_15_local_g0_3_69868)
  );
  LocalMux t6005 (
    .I(seg_14_14_sp4_h_r_20_54525),
    .O(seg_14_14_local_g0_4_58254)
  );
  Span4Mux_h3 t6006 (
    .I(seg_17_14_sp4_v_t_38_66142),
    .O(seg_14_14_sp4_h_r_20_54525)
  );
  LocalMux t6007 (
    .I(seg_17_10_sp4_h_r_4_69350),
    .O(seg_17_10_local_g0_4_69254)
  );
  Span4Mux_h0 t6008 (
    .I(seg_17_10_sp4_v_t_46_65658),
    .O(seg_17_10_sp4_h_r_4_69350)
  );
  Span4Mux_v4 t6009 (
    .I(seg_17_14_sp4_v_t_38_66142),
    .O(seg_17_10_sp4_v_t_46_65658)
  );
  CascadeMux t601 (
    .I(net_45446),
    .O(net_45446_cascademuxed)
  );
  LocalMux t6010 (
    .I(seg_16_17_neigh_op_tnr_6_66368),
    .O(seg_16_17_local_g2_6_66302)
  );
  LocalMux t6011 (
    .I(seg_17_17_neigh_op_top_6_66368),
    .O(seg_17_17_local_g0_6_70117)
  );
  LocalMux t6012 (
    .I(seg_14_18_sp4_h_r_9_58847),
    .O(seg_14_18_local_g1_1_58751)
  );
  LocalMux t6013 (
    .I(seg_16_16_sp4_r_v_b_7_65900),
    .O(seg_16_16_local_g1_7_66172)
  );
  Span4Mux_v1 t6014 (
    .I(seg_17_16_sp4_v_t_41_66391),
    .O(seg_16_16_sp4_r_v_b_7_65900)
  );
  LocalMux t6015 (
    .I(seg_17_14_sp4_v_b_31_65900),
    .O(seg_17_14_local_g2_7_69765)
  );
  Span4Mux_v2 t6016 (
    .I(seg_17_16_sp4_v_t_41_66391),
    .O(seg_17_14_sp4_v_b_31_65900)
  );
  LocalMux t6017 (
    .I(seg_17_14_sp4_v_b_31_65900),
    .O(seg_17_14_local_g3_7_69773)
  );
  LocalMux t6018 (
    .I(seg_4_3_sp4_h_r_16_15489),
    .O(seg_4_3_local_g0_0_19219)
  );
  Span4Mux_h3 t6019 (
    .I(seg_7_3_sp4_h_r_9_30186),
    .O(seg_4_3_sp4_h_r_16_15489)
  );
  CascadeMux t602 (
    .I(net_45452),
    .O(net_45452_cascademuxed)
  );
  Span4Mux_h4 t6020 (
    .I(seg_11_3_sp4_h_r_6_45507),
    .O(seg_7_3_sp4_h_r_9_30186)
  );
  Span4Mux_h4 t6021 (
    .I(seg_15_3_sp4_v_b_1_56739),
    .O(seg_11_3_sp4_h_r_6_45507)
  );
  IoSpan4Mux t6022 (
    .I(seg_15_0_span4_horz_r_0_60431),
    .O(seg_15_3_sp4_v_b_1_56739)
  );
  LocalMux t6023 (
    .I(seg_4_3_sp4_h_r_15_15486),
    .O(seg_4_3_local_g1_7_19234)
  );
  Span4Mux_h3 t6024 (
    .I(seg_7_3_sp4_h_r_6_30183),
    .O(seg_4_3_sp4_h_r_15_15486)
  );
  Span4Mux_h4 t6025 (
    .I(seg_11_3_sp4_h_r_6_45507),
    .O(seg_7_3_sp4_h_r_6_30183)
  );
  LocalMux t6026 (
    .I(seg_16_3_sp4_v_b_43_60840),
    .O(seg_16_3_local_g3_3_64585)
  );
  Span4Mux_v1 t6027 (
    .I(seg_16_2_sp4_h_r_0_64529),
    .O(seg_16_3_sp4_v_b_43_60840)
  );
  LocalMux t6028 (
    .I(seg_7_0_span4_vert_15_26690),
    .O(seg_7_0_local_g1_7_29752)
  );
  Span4Mux_v2 t6029 (
    .I(seg_7_2_sp4_h_r_9_30063),
    .O(seg_7_0_span4_vert_15_26690)
  );
  CascadeMux t603 (
    .I(net_45458),
    .O(net_45458_cascademuxed)
  );
  Span4Mux_h4 t6030 (
    .I(seg_11_2_sp4_h_r_1_45377),
    .O(seg_7_2_sp4_h_r_9_30063)
  );
  Span4Mux_h4 t6031 (
    .I(seg_15_2_sp4_h_r_5_60705),
    .O(seg_11_2_sp4_h_r_1_45377)
  );
  LocalMux t6032 (
    .I(seg_18_4_neigh_op_bot_0_68348),
    .O(seg_18_4_local_g1_0_72351)
  );
  LocalMux t6033 (
    .I(seg_18_4_neigh_op_bot_1_68349),
    .O(seg_18_4_local_g0_1_72344)
  );
  LocalMux t6034 (
    .I(seg_18_4_neigh_op_bot_2_68350),
    .O(seg_18_4_local_g1_2_72353)
  );
  LocalMux t6035 (
    .I(seg_18_4_neigh_op_bot_3_68351),
    .O(seg_18_4_local_g0_3_72346)
  );
  LocalMux t6036 (
    .I(seg_18_4_neigh_op_bot_4_68352),
    .O(seg_18_4_local_g1_4_72355)
  );
  LocalMux t6037 (
    .I(seg_18_3_lutff_5_out_68353),
    .O(seg_18_3_local_g3_5_72249)
  );
  LocalMux t6038 (
    .I(seg_18_4_neigh_op_bot_7_68355),
    .O(seg_18_4_local_g1_7_72358)
  );
  LocalMux t6039 (
    .I(seg_18_5_sp4_v_b_20_68503),
    .O(seg_18_5_local_g1_4_72478)
  );
  CascadeMux t604 (
    .I(net_45464),
    .O(net_45464_cascademuxed)
  );
  LocalMux t6040 (
    .I(seg_18_7_sp4_v_b_21_68750),
    .O(seg_18_7_local_g0_5_72717)
  );
  Span4Mux_v3 t6041 (
    .I(seg_18_4_sp4_h_r_2_72441),
    .O(seg_18_7_sp4_v_b_21_68750)
  );
  LocalMux t6042 (
    .I(seg_18_7_sp4_r_v_b_8_72458),
    .O(seg_18_7_local_g2_0_72728)
  );
  LocalMux t6043 (
    .I(seg_18_7_sp4_r_v_b_10_72460),
    .O(seg_18_7_local_g2_2_72730)
  );
  LocalMux t6044 (
    .I(seg_18_7_sp4_v_b_1_68618),
    .O(seg_18_7_local_g1_1_72721)
  );
  LocalMux t6045 (
    .I(seg_18_7_sp4_v_b_3_68620),
    .O(seg_18_7_local_g1_3_72723)
  );
  LocalMux t6046 (
    .I(seg_18_7_sp4_v_b_5_68622),
    .O(seg_18_7_local_g1_5_72725)
  );
  LocalMux t6047 (
    .I(seg_18_7_sp4_v_b_7_68624),
    .O(seg_18_7_local_g1_7_72727)
  );
  LocalMux t6048 (
    .I(seg_18_4_neigh_op_top_2_68596),
    .O(seg_18_4_local_g0_2_72345)
  );
  LocalMux t6049 (
    .I(seg_18_6_neigh_op_bot_2_68596),
    .O(seg_18_6_local_g1_2_72599)
  );
  CascadeMux t605 (
    .I(net_45470),
    .O(net_45470_cascademuxed)
  );
  LocalMux t6050 (
    .I(seg_18_5_lutff_3_out_68597),
    .O(seg_18_5_local_g0_3_72469)
  );
  LocalMux t6051 (
    .I(seg_18_4_neigh_op_top_4_68598),
    .O(seg_18_4_local_g0_4_72347)
  );
  LocalMux t6052 (
    .I(seg_18_5_lutff_5_out_68599),
    .O(seg_18_5_local_g3_5_72495)
  );
  LocalMux t6053 (
    .I(seg_18_4_neigh_op_top_6_68600),
    .O(seg_18_4_local_g0_6_72349)
  );
  LocalMux t6054 (
    .I(seg_18_4_neigh_op_top_7_68601),
    .O(seg_18_4_local_g0_7_72350)
  );
  LocalMux t6055 (
    .I(seg_18_8_sp4_v_b_19_68871),
    .O(seg_18_8_local_g1_3_72846)
  );
  Span4Mux_v3 t6056 (
    .I(seg_18_5_sp4_h_r_0_72560),
    .O(seg_18_8_sp4_v_b_19_68871)
  );
  LocalMux t6057 (
    .I(seg_18_8_sp4_v_b_15_68867),
    .O(seg_18_8_local_g1_7_72850)
  );
  Span4Mux_v3 t6058 (
    .I(seg_18_5_sp4_h_r_2_72564),
    .O(seg_18_8_sp4_v_b_15_68867)
  );
  LocalMux t6059 (
    .I(seg_18_6_lutff_1_out_68718),
    .O(seg_18_6_local_g0_1_72590)
  );
  CascadeMux t606 (
    .I(net_45476),
    .O(net_45476_cascademuxed)
  );
  LocalMux t6060 (
    .I(seg_17_6_neigh_op_rgt_3_68720),
    .O(seg_17_6_local_g3_3_68785)
  );
  LocalMux t6061 (
    .I(seg_18_5_neigh_op_top_5_68722),
    .O(seg_18_5_local_g1_5_72479)
  );
  LocalMux t6062 (
    .I(seg_18_5_neigh_op_top_6_68723),
    .O(seg_18_5_local_g0_6_72472)
  );
  LocalMux t6063 (
    .I(seg_18_7_neigh_op_bot_7_68724),
    .O(seg_18_7_local_g0_7_72719)
  );
  LocalMux t6064 (
    .I(seg_16_7_sp4_h_r_15_61317),
    .O(seg_16_7_local_g1_7_65065)
  );
  Span4Mux_h3 t6065 (
    .I(seg_19_7_sp4_v_b_2_72452),
    .O(seg_16_7_sp4_h_r_15_61317)
  );
  LocalMux t6066 (
    .I(seg_18_4_sp4_v_b_24_68496),
    .O(seg_18_4_local_g2_0_72359)
  );
  LocalMux t6067 (
    .I(seg_17_4_sp4_r_v_b_32_68504),
    .O(seg_17_4_local_g0_3_68515)
  );
  LocalMux t6068 (
    .I(seg_11_17_sp12_v_b_5_45989),
    .O(seg_11_17_local_g3_5_47156)
  );
  Span12Mux_v10 t6069 (
    .I(seg_11_7_sp12_h_r_1_45988),
    .O(seg_11_17_sp12_v_b_5_45989)
  );
  CascadeMux t607 (
    .I(net_45563),
    .O(net_45563_cascademuxed)
  );
  LocalMux t6070 (
    .I(seg_10_16_sp12_v_b_7_42159),
    .O(seg_10_16_local_g2_7_43196)
  );
  Span12Mux_v9 t6071 (
    .I(seg_10_7_sp12_h_r_0_42156),
    .O(seg_10_16_sp12_v_b_7_42159)
  );
  LocalMux t6072 (
    .I(seg_9_15_sp12_v_b_9_38327),
    .O(seg_9_15_local_g2_1_39236)
  );
  Span12Mux_v8 t6073 (
    .I(seg_9_7_sp12_h_r_1_38326),
    .O(seg_9_15_sp12_v_b_9_38327)
  );
  LocalMux t6074 (
    .I(seg_9_16_sp12_h_r_6_28234),
    .O(seg_9_16_local_g0_6_39348)
  );
  Span12Mux_h9 t6075 (
    .I(seg_18_16_sp12_v_b_1_72435),
    .O(seg_9_16_sp12_h_r_6_28234)
  );
  LocalMux t6076 (
    .I(seg_10_16_sp12_h_r_9_28234),
    .O(seg_10_16_local_g1_1_43182)
  );
  Span12Mux_h8 t6077 (
    .I(seg_18_16_sp12_v_b_1_72435),
    .O(seg_10_16_sp12_h_r_9_28234)
  );
  LocalMux t6078 (
    .I(seg_13_14_sp4_v_b_21_50458),
    .O(seg_13_14_local_g0_5_54425)
  );
  Span4Mux_v3 t6079 (
    .I(seg_13_11_sp4_h_r_2_54149),
    .O(seg_13_14_sp4_v_b_21_50458)
  );
  CascadeMux t608 (
    .I(net_45569),
    .O(net_45569_cascademuxed)
  );
  Span4Mux_h4 t6080 (
    .I(seg_17_11_sp4_v_b_9_65287),
    .O(seg_13_11_sp4_h_r_2_54149)
  );
  Span4Mux_v4 t6081 (
    .I(seg_17_7_sp4_h_r_3_68980),
    .O(seg_17_11_sp4_v_b_9_65287)
  );
  LocalMux t6082 (
    .I(seg_13_15_sp4_v_b_8_50458),
    .O(seg_13_15_local_g0_0_54543)
  );
  Span4Mux_v4 t6083 (
    .I(seg_13_11_sp4_h_r_2_54149),
    .O(seg_13_15_sp4_v_b_8_50458)
  );
  LocalMux t6084 (
    .I(seg_20_14_sp4_r_v_b_19_80471),
    .O(seg_20_14_local_g3_3_80631)
  );
  Span4Mux_v3 t6085 (
    .I(seg_21_11_sp4_v_b_3_79974),
    .O(seg_20_14_sp4_r_v_b_19_80471)
  );
  Span4Mux_v4 t6086 (
    .I(seg_21_7_sp4_h_l_38_68980),
    .O(seg_21_11_sp4_v_b_3_79974)
  );
  LocalMux t6087 (
    .I(seg_10_14_sp4_v_b_16_38960),
    .O(seg_10_14_local_g0_0_42927)
  );
  Span4Mux_v3 t6088 (
    .I(seg_10_11_sp4_v_b_5_38468),
    .O(seg_10_14_sp4_v_b_16_38960)
  );
  Span4Mux_v4 t6089 (
    .I(seg_10_7_sp4_h_r_5_42167),
    .O(seg_10_11_sp4_v_b_5_38468)
  );
  CascadeMux t609 (
    .I(net_45575),
    .O(net_45575_cascademuxed)
  );
  Span4Mux_h4 t6090 (
    .I(seg_14_7_sp4_h_r_5_57490),
    .O(seg_10_7_sp4_h_r_5_42167)
  );
  Span4Mux_h4 t6091 (
    .I(seg_18_7_sp4_h_r_2_72810),
    .O(seg_14_7_sp4_h_r_5_57490)
  );
  LocalMux t6092 (
    .I(seg_13_15_sp4_h_r_8_54647),
    .O(seg_13_15_local_g1_0_54551)
  );
  Span4Mux_h4 t6093 (
    .I(seg_17_15_sp4_v_b_3_65773),
    .O(seg_13_15_sp4_h_r_8_54647)
  );
  Span4Mux_v4 t6094 (
    .I(seg_17_11_sp4_v_b_3_65281),
    .O(seg_17_15_sp4_v_b_3_65773)
  );
  Span4Mux_v4 t6095 (
    .I(seg_17_7_sp4_h_r_9_68986),
    .O(seg_17_11_sp4_v_b_3_65281)
  );
  LocalMux t6096 (
    .I(seg_13_15_sp4_h_r_18_50815),
    .O(seg_13_15_local_g1_2_54553)
  );
  Span4Mux_h3 t6097 (
    .I(seg_16_15_sp4_v_b_7_61946),
    .O(seg_13_15_sp4_h_r_18_50815)
  );
  Span4Mux_v4 t6098 (
    .I(seg_16_11_sp4_v_b_4_61453),
    .O(seg_16_15_sp4_v_b_7_61946)
  );
  Span4Mux_v4 t6099 (
    .I(seg_16_7_sp4_h_r_4_65150),
    .O(seg_16_11_sp4_v_b_4_61453)
  );
  CascadeMux t61 (
    .I(net_11469),
    .O(net_11469_cascademuxed)
  );
  CascadeMux t610 (
    .I(net_45581),
    .O(net_45581_cascademuxed)
  );
  LocalMux t6100 (
    .I(seg_10_14_sp4_r_v_b_17_42792),
    .O(seg_10_14_local_g3_1_42952)
  );
  Span4Mux_v3 t6101 (
    .I(seg_11_11_sp4_v_b_1_42295),
    .O(seg_10_14_sp4_r_v_b_17_42792)
  );
  Span4Mux_v4 t6102 (
    .I(seg_11_7_sp4_h_r_1_45992),
    .O(seg_11_11_sp4_v_b_1_42295)
  );
  Span4Mux_h4 t6103 (
    .I(seg_15_7_sp4_h_r_5_61320),
    .O(seg_11_7_sp4_h_r_1_45992)
  );
  LocalMux t6104 (
    .I(seg_11_15_sp4_v_b_7_42793),
    .O(seg_11_15_local_g1_7_46896)
  );
  Span4Mux_v4 t6105 (
    .I(seg_11_11_sp4_h_r_7_46492),
    .O(seg_11_15_sp4_v_b_7_42793)
  );
  Span4Mux_h4 t6106 (
    .I(seg_15_11_sp4_v_b_7_57624),
    .O(seg_11_11_sp4_h_r_7_46492)
  );
  Span4Mux_v4 t6107 (
    .I(seg_15_7_sp4_h_r_7_61322),
    .O(seg_15_11_sp4_v_b_7_57624)
  );
  LocalMux t6108 (
    .I(seg_13_12_sp4_r_v_b_2_53914),
    .O(seg_13_12_local_g1_2_54184)
  );
  Span4Mux_v4 t6109 (
    .I(seg_14_8_sp4_h_r_8_57616),
    .O(seg_13_12_sp4_r_v_b_2_53914)
  );
  CascadeMux t611 (
    .I(net_45587),
    .O(net_45587_cascademuxed)
  );
  Span4Mux_h4 t6110 (
    .I(seg_18_8_sp4_v_b_3_68743),
    .O(seg_14_8_sp4_h_r_8_57616)
  );
  LocalMux t6111 (
    .I(seg_9_16_sp4_r_v_b_14_39204),
    .O(seg_9_16_local_g2_6_39364)
  );
  Span4Mux_v3 t6112 (
    .I(seg_10_13_sp4_h_r_9_42909),
    .O(seg_9_16_sp4_r_v_b_14_39204)
  );
  Span4Mux_h4 t6113 (
    .I(seg_14_13_sp4_h_r_1_58222),
    .O(seg_10_13_sp4_h_r_9_42909)
  );
  Span4Mux_h4 t6114 (
    .I(seg_18_13_sp4_v_b_8_69365),
    .O(seg_14_13_sp4_h_r_1_58222)
  );
  Span4Mux_v4 t6115 (
    .I(seg_18_9_sp4_v_b_0_68865),
    .O(seg_18_13_sp4_v_b_8_69365)
  );
  LocalMux t6116 (
    .I(seg_11_17_sp4_h_r_12_43391),
    .O(seg_11_17_local_g0_4_47131)
  );
  Span4Mux_h3 t6117 (
    .I(seg_14_17_sp4_v_b_1_54526),
    .O(seg_11_17_sp4_h_r_12_43391)
  );
  Span4Mux_v4 t6118 (
    .I(seg_14_13_sp4_h_r_1_58222),
    .O(seg_14_17_sp4_v_b_1_54526)
  );
  LocalMux t6119 (
    .I(seg_13_12_sp4_r_v_b_14_54036),
    .O(seg_13_12_local_g2_6_54196)
  );
  CascadeMux t612 (
    .I(net_45593),
    .O(net_45593_cascademuxed)
  );
  Span4Mux_v3 t6120 (
    .I(seg_14_9_sp4_h_r_9_57740),
    .O(seg_13_12_sp4_r_v_b_14_54036)
  );
  Span4Mux_h4 t6121 (
    .I(seg_18_9_sp4_v_b_4_68869),
    .O(seg_14_9_sp4_h_r_9_57740)
  );
  LocalMux t6122 (
    .I(seg_9_17_sp4_r_v_b_9_39210),
    .O(seg_9_17_local_g2_1_39482)
  );
  Span4Mux_v4 t6123 (
    .I(seg_10_13_sp4_v_b_9_38718),
    .O(seg_9_17_sp4_r_v_b_9_39210)
  );
  Span4Mux_v4 t6124 (
    .I(seg_10_9_sp4_h_r_3_42411),
    .O(seg_10_13_sp4_v_b_9_38718)
  );
  Span4Mux_h4 t6125 (
    .I(seg_14_9_sp4_h_r_3_57734),
    .O(seg_10_9_sp4_h_r_3_42411)
  );
  Span4Mux_h4 t6126 (
    .I(seg_18_9_sp4_v_b_10_68875),
    .O(seg_14_9_sp4_h_r_3_57734)
  );
  LocalMux t6127 (
    .I(seg_13_12_sp4_r_v_b_25_54157),
    .O(seg_13_12_local_g1_1_54183)
  );
  Span4Mux_v2 t6128 (
    .I(seg_14_10_sp4_h_r_1_57853),
    .O(seg_13_12_sp4_r_v_b_25_54157)
  );
  Span4Mux_h4 t6129 (
    .I(seg_18_10_sp4_v_b_1_68987),
    .O(seg_14_10_sp4_h_r_1_57853)
  );
  CascadeMux t613 (
    .I(net_45599),
    .O(net_45599_cascademuxed)
  );
  LocalMux t6130 (
    .I(seg_13_13_sp4_r_v_b_12_54157),
    .O(seg_13_13_local_g2_4_54317)
  );
  Span4Mux_v3 t6131 (
    .I(seg_14_10_sp4_h_r_1_57853),
    .O(seg_13_13_sp4_r_v_b_12_54157)
  );
  LocalMux t6132 (
    .I(seg_13_14_sp4_r_v_b_1_54157),
    .O(seg_13_14_local_g1_1_54429)
  );
  Span4Mux_v4 t6133 (
    .I(seg_14_10_sp4_h_r_1_57853),
    .O(seg_13_14_sp4_r_v_b_1_54157)
  );
  LocalMux t6134 (
    .I(seg_9_16_sp4_r_v_b_27_39327),
    .O(seg_9_16_local_g0_3_39345)
  );
  Span4Mux_v2 t6135 (
    .I(seg_10_14_sp4_h_r_3_43026),
    .O(seg_9_16_sp4_r_v_b_27_39327)
  );
  Span4Mux_h4 t6136 (
    .I(seg_14_14_sp4_h_r_3_58349),
    .O(seg_10_14_sp4_h_r_3_43026)
  );
  Span4Mux_h4 t6137 (
    .I(seg_18_14_sp4_v_b_3_69481),
    .O(seg_14_14_sp4_h_r_3_58349)
  );
  Span4Mux_v4 t6138 (
    .I(seg_18_10_sp4_v_b_3_68989),
    .O(seg_18_14_sp4_v_b_3_69481)
  );
  LocalMux t6139 (
    .I(seg_10_16_sp4_v_b_27_39327),
    .O(seg_10_16_local_g2_3_43192)
  );
  CascadeMux t614 (
    .I(net_45605),
    .O(net_45605_cascademuxed)
  );
  Span4Mux_v2 t6140 (
    .I(seg_10_14_sp4_h_r_3_43026),
    .O(seg_10_16_sp4_v_b_27_39327)
  );
  LocalMux t6141 (
    .I(seg_10_17_sp4_v_b_14_39327),
    .O(seg_10_17_local_g1_6_43310)
  );
  Span4Mux_v3 t6142 (
    .I(seg_10_14_sp4_h_r_3_43026),
    .O(seg_10_17_sp4_v_b_14_39327)
  );
  LocalMux t6143 (
    .I(seg_10_14_sp4_v_b_9_38841),
    .O(seg_10_14_local_g1_1_42936)
  );
  Span4Mux_v4 t6144 (
    .I(seg_10_10_sp4_h_r_3_42534),
    .O(seg_10_14_sp4_v_b_9_38841)
  );
  Span4Mux_h4 t6145 (
    .I(seg_14_10_sp4_h_r_0_57852),
    .O(seg_10_10_sp4_h_r_3_42534)
  );
  Span4Mux_h4 t6146 (
    .I(seg_18_10_sp4_v_b_7_68993),
    .O(seg_14_10_sp4_h_r_0_57852)
  );
  LocalMux t6147 (
    .I(seg_13_12_sp4_r_v_b_30_54164),
    .O(seg_13_12_local_g0_6_54180)
  );
  Span4Mux_v2 t6148 (
    .I(seg_14_10_sp4_h_r_0_57852),
    .O(seg_13_12_sp4_r_v_b_30_54164)
  );
  LocalMux t6149 (
    .I(seg_13_13_sp4_r_v_b_20_54165),
    .O(seg_13_13_local_g3_4_54325)
  );
  CascadeMux t615 (
    .I(net_45692),
    .O(net_45692_cascademuxed)
  );
  Span4Mux_v3 t6150 (
    .I(seg_14_10_sp4_h_r_9_57863),
    .O(seg_13_13_sp4_r_v_b_20_54165)
  );
  Span4Mux_h4 t6151 (
    .I(seg_18_10_sp4_v_b_9_68995),
    .O(seg_14_10_sp4_h_r_9_57863)
  );
  LocalMux t6152 (
    .I(seg_13_14_sp4_r_v_b_9_54165),
    .O(seg_13_14_local_g2_1_54437)
  );
  Span4Mux_v4 t6153 (
    .I(seg_14_10_sp4_h_r_9_57863),
    .O(seg_13_14_sp4_r_v_b_9_54165)
  );
  LocalMux t6154 (
    .I(seg_13_15_sp4_r_v_b_16_54407),
    .O(seg_13_15_local_g3_0_54567)
  );
  Span4Mux_v3 t6155 (
    .I(seg_14_12_sp4_h_r_11_58101),
    .O(seg_13_15_sp4_r_v_b_16_54407)
  );
  Span4Mux_h4 t6156 (
    .I(seg_18_12_sp4_v_b_6_69240),
    .O(seg_14_12_sp4_h_r_11_58101)
  );
  Span4Mux_v4 t6157 (
    .I(seg_18_8_sp4_h_r_0_72929),
    .O(seg_18_12_sp4_v_b_6_69240)
  );
  LocalMux t6158 (
    .I(seg_13_7_sp4_v_b_13_49589),
    .O(seg_13_7_local_g0_5_53564)
  );
  Span4Mux_v1 t6159 (
    .I(seg_13_8_sp4_h_r_7_53785),
    .O(seg_13_7_sp4_v_b_13_49589)
  );
  CascadeMux t616 (
    .I(net_46055),
    .O(net_46055_cascademuxed)
  );
  Span4Mux_h4 t6160 (
    .I(seg_17_8_sp4_h_r_7_69107),
    .O(seg_13_8_sp4_h_r_7_53785)
  );
  LocalMux t6161 (
    .I(seg_13_10_sp4_r_v_b_34_53922),
    .O(seg_13_10_local_g0_1_53929)
  );
  Span4Mux_v2 t6162 (
    .I(seg_14_8_sp4_h_r_10_57608),
    .O(seg_13_10_sp4_r_v_b_34_53922)
  );
  Span4Mux_h4 t6163 (
    .I(seg_18_8_sp4_h_r_2_72933),
    .O(seg_14_8_sp4_h_r_10_57608)
  );
  LocalMux t6164 (
    .I(seg_14_11_sp4_v_b_23_53922),
    .O(seg_14_11_local_g1_7_57896)
  );
  Span4Mux_v3 t6165 (
    .I(seg_14_8_sp4_h_r_10_57608),
    .O(seg_14_11_sp4_v_b_23_53922)
  );
  LocalMux t6166 (
    .I(seg_11_15_sp4_r_v_b_13_46742),
    .O(seg_11_15_local_g2_5_46902)
  );
  Span4Mux_v3 t6167 (
    .I(seg_12_12_sp4_v_b_4_46254),
    .O(seg_11_15_sp4_r_v_b_13_46742)
  );
  Span4Mux_v4 t6168 (
    .I(seg_12_8_sp4_h_r_4_49951),
    .O(seg_12_12_sp4_v_b_4_46254)
  );
  Span4Mux_h4 t6169 (
    .I(seg_16_8_sp4_h_r_8_65277),
    .O(seg_12_8_sp4_h_r_4_49951)
  );
  CascadeMux t617 (
    .I(net_46061),
    .O(net_46061_cascademuxed)
  );
  LocalMux t6170 (
    .I(seg_15_8_sp4_h_r_5_61443),
    .O(seg_15_8_local_g0_5_61347)
  );
  LocalMux t6171 (
    .I(seg_15_8_sp4_h_r_11_61439),
    .O(seg_15_8_local_g0_3_61345)
  );
  LocalMux t6172 (
    .I(seg_15_9_sp4_h_r_11_61562),
    .O(seg_15_9_local_g0_3_61468)
  );
  Span4Mux_h4 t6173 (
    .I(seg_19_9_sp4_v_b_6_72702),
    .O(seg_15_9_sp4_h_r_11_61562)
  );
  LocalMux t6174 (
    .I(seg_17_5_sp4_r_v_b_47_68752),
    .O(seg_17_5_local_g3_7_68666)
  );
  LocalMux t6175 (
    .I(seg_9_14_sp4_r_v_b_10_38844),
    .O(seg_9_14_local_g2_2_39114)
  );
  Span4Mux_v4 t6176 (
    .I(seg_10_10_sp4_h_r_4_42535),
    .O(seg_9_14_sp4_r_v_b_10_38844)
  );
  Span4Mux_h4 t6177 (
    .I(seg_14_10_sp4_h_r_8_57862),
    .O(seg_10_10_sp4_h_r_4_42535)
  );
  Span4Mux_h4 t6178 (
    .I(seg_18_10_sp4_v_b_8_68996),
    .O(seg_14_10_sp4_h_r_8_57862)
  );
  LocalMux t6179 (
    .I(seg_13_14_sp4_r_v_b_8_54166),
    .O(seg_13_14_local_g2_0_54436)
  );
  CascadeMux t618 (
    .I(net_46079),
    .O(net_46079_cascademuxed)
  );
  Span4Mux_v4 t6180 (
    .I(seg_14_10_sp4_h_r_8_57862),
    .O(seg_13_14_sp4_r_v_b_8_54166)
  );
  LocalMux t6181 (
    .I(seg_18_9_lutff_0_out_69086),
    .O(seg_18_9_local_g2_0_72974)
  );
  LocalMux t6182 (
    .I(seg_18_9_lutff_5_out_69091),
    .O(seg_18_9_local_g3_5_72987)
  );
  LocalMux t6183 (
    .I(seg_18_10_neigh_op_bot_5_69091),
    .O(seg_18_10_local_g1_5_73094)
  );
  LocalMux t6184 (
    .I(seg_18_10_neigh_op_bot_6_69092),
    .O(seg_18_10_local_g0_6_73087)
  );
  LocalMux t6185 (
    .I(seg_20_4_sp4_v_b_13_75992),
    .O(seg_20_4_local_g1_5_79387)
  );
  Span4Mux_v1 t6186 (
    .I(seg_20_5_sp4_v_t_41_76404),
    .O(seg_20_4_sp4_v_b_13_75992)
  );
  Span4Mux_v4 t6187 (
    .I(seg_20_9_sp4_h_l_47_65392),
    .O(seg_20_5_sp4_v_t_41_76404)
  );
  LocalMux t6188 (
    .I(seg_20_10_sp4_h_r_23_76797),
    .O(seg_20_10_local_g1_7_80127)
  );
  Span4Mux_h1 t6189 (
    .I(seg_19_10_sp4_v_b_10_72829),
    .O(seg_20_10_sp4_h_r_23_76797)
  );
  CascadeMux t619 (
    .I(net_46307),
    .O(net_46307_cascademuxed)
  );
  LocalMux t6190 (
    .I(seg_18_10_lutff_1_out_69210),
    .O(seg_18_10_local_g3_1_73106)
  );
  LocalMux t6191 (
    .I(seg_17_10_neigh_op_rgt_3_69212),
    .O(seg_17_10_local_g2_3_69269)
  );
  LocalMux t6192 (
    .I(seg_18_9_neigh_op_top_4_69213),
    .O(seg_18_9_local_g1_4_72970)
  );
  LocalMux t6193 (
    .I(seg_17_10_neigh_op_rgt_6_69215),
    .O(seg_17_10_local_g3_6_69280)
  );
  LocalMux t6194 (
    .I(seg_20_9_sp4_v_b_15_76504),
    .O(seg_20_9_local_g0_7_79996)
  );
  Span4Mux_v1 t6195 (
    .I(seg_20_10_sp4_h_l_39_65517),
    .O(seg_20_9_sp4_v_b_15_76504)
  );
  LocalMux t6196 (
    .I(seg_20_10_sp4_h_r_6_80214),
    .O(seg_20_10_local_g0_6_80118)
  );
  Span4Mux_h0 t6197 (
    .I(seg_20_10_sp4_h_l_43_65521),
    .O(seg_20_10_sp4_h_r_6_80214)
  );
  LocalMux t6198 (
    .I(seg_20_11_sp4_h_r_15_76901),
    .O(seg_20_11_local_g0_7_80242)
  );
  Span4Mux_h1 t6199 (
    .I(seg_19_11_sp4_v_b_8_72950),
    .O(seg_20_11_sp4_h_r_15_76901)
  );
  CascadeMux t62 (
    .I(net_11475),
    .O(net_11475_cascademuxed)
  );
  CascadeMux t620 (
    .I(net_46343),
    .O(net_46343_cascademuxed)
  );
  LocalMux t6200 (
    .I(seg_17_11_neigh_op_rgt_0_69332),
    .O(seg_17_11_local_g3_0_69397)
  );
  LocalMux t6201 (
    .I(seg_18_11_lutff_1_out_69333),
    .O(seg_18_11_local_g0_1_73205)
  );
  LocalMux t6202 (
    .I(seg_17_11_neigh_op_rgt_2_69334),
    .O(seg_17_11_local_g3_2_69399)
  );
  LocalMux t6203 (
    .I(seg_18_11_lutff_3_out_69335),
    .O(seg_18_11_local_g2_3_73223)
  );
  LocalMux t6204 (
    .I(seg_18_11_lutff_5_out_69337),
    .O(seg_18_11_local_g2_5_73225)
  );
  LocalMux t6205 (
    .I(seg_18_11_lutff_6_out_69338),
    .O(seg_18_11_local_g1_6_73218)
  );
  LocalMux t6206 (
    .I(seg_18_10_neigh_op_top_7_69339),
    .O(seg_18_10_local_g1_7_73096)
  );
  LocalMux t6207 (
    .I(seg_12_12_sp4_v_b_44_46626),
    .O(seg_12_12_local_g2_4_50363)
  );
  Span4Mux_v1 t6208 (
    .I(seg_12_11_sp4_h_r_3_50319),
    .O(seg_12_12_sp4_v_b_44_46626)
  );
  Span4Mux_h4 t6209 (
    .I(seg_16_11_sp4_h_r_0_65636),
    .O(seg_12_11_sp4_h_r_3_50319)
  );
  CascadeMux t621 (
    .I(net_46424),
    .O(net_46424_cascademuxed)
  );
  LocalMux t6210 (
    .I(seg_12_11_sp4_h_r_21_46493),
    .O(seg_12_11_local_g1_5_50233)
  );
  Span4Mux_h3 t6211 (
    .I(seg_15_11_sp4_h_r_5_61812),
    .O(seg_12_11_sp4_h_r_21_46493)
  );
  LocalMux t6212 (
    .I(seg_14_11_sp4_h_r_4_57981),
    .O(seg_14_11_local_g1_4_57893)
  );
  Span4Mux_h4 t6213 (
    .I(seg_18_11_sp4_h_r_8_73308),
    .O(seg_14_11_sp4_h_r_4_57981)
  );
  LocalMux t6214 (
    .I(seg_13_12_sp4_r_v_b_23_54045),
    .O(seg_13_12_local_g3_7_54205)
  );
  Span4Mux_v1 t6215 (
    .I(seg_14_13_sp4_h_r_5_58228),
    .O(seg_13_12_sp4_r_v_b_23_54045)
  );
  Span4Mux_h4 t6216 (
    .I(seg_18_13_sp4_v_b_0_69357),
    .O(seg_14_13_sp4_h_r_5_58228)
  );
  LocalMux t6217 (
    .I(seg_17_11_neigh_op_tnr_0_69455),
    .O(seg_17_11_local_g2_0_69389)
  );
  LocalMux t6218 (
    .I(seg_18_12_lutff_1_out_69456),
    .O(seg_18_12_local_g3_1_73352)
  );
  LocalMux t6219 (
    .I(seg_17_11_neigh_op_tnr_2_69457),
    .O(seg_17_11_local_g2_2_69391)
  );
  CascadeMux t622 (
    .I(net_46442),
    .O(net_46442_cascademuxed)
  );
  LocalMux t6220 (
    .I(seg_18_12_lutff_3_out_69458),
    .O(seg_18_12_local_g0_3_73330)
  );
  LocalMux t6221 (
    .I(seg_18_12_lutff_4_out_69459),
    .O(seg_18_12_local_g0_4_73331)
  );
  LocalMux t6222 (
    .I(seg_17_11_neigh_op_tnr_6_69461),
    .O(seg_17_11_local_g3_6_69403)
  );
  LocalMux t6223 (
    .I(seg_18_10_sp4_v_b_38_69358),
    .O(seg_18_10_local_g2_6_73103)
  );
  LocalMux t6224 (
    .I(seg_18_12_neigh_op_top_0_69578),
    .O(seg_18_12_local_g1_0_73335)
  );
  LocalMux t6225 (
    .I(seg_16_13_sp4_h_r_10_65884),
    .O(seg_16_13_local_g0_2_65790)
  );
  LocalMux t6226 (
    .I(seg_16_13_sp4_h_r_12_62052),
    .O(seg_16_13_local_g0_4_65792)
  );
  LocalMux t6227 (
    .I(seg_16_13_sp4_h_r_16_62058),
    .O(seg_16_13_local_g1_0_65796)
  );
  LocalMux t6228 (
    .I(seg_16_13_sp4_h_r_20_62062),
    .O(seg_16_13_local_g1_4_65800)
  );
  LocalMux t6229 (
    .I(seg_18_10_sp4_v_b_47_69367),
    .O(seg_18_10_local_g2_7_73104)
  );
  CascadeMux t623 (
    .I(net_46547),
    .O(net_46547_cascademuxed)
  );
  LocalMux t6230 (
    .I(seg_18_15_neigh_op_bot_0_69701),
    .O(seg_18_15_local_g1_0_73704)
  );
  LocalMux t6231 (
    .I(seg_18_13_neigh_op_top_1_69702),
    .O(seg_18_13_local_g1_1_73459)
  );
  LocalMux t6232 (
    .I(seg_18_15_neigh_op_bot_2_69703),
    .O(seg_18_15_local_g0_2_73698)
  );
  LocalMux t6233 (
    .I(seg_18_15_neigh_op_bot_3_69704),
    .O(seg_18_15_local_g1_3_73707)
  );
  LocalMux t6234 (
    .I(seg_18_15_neigh_op_bot_4_69705),
    .O(seg_18_15_local_g1_4_73708)
  );
  LocalMux t6235 (
    .I(seg_18_15_neigh_op_bot_7_69708),
    .O(seg_18_15_local_g1_7_73711)
  );
  LocalMux t6236 (
    .I(seg_16_14_sp4_h_r_6_66013),
    .O(seg_16_14_local_g0_6_65917)
  );
  LocalMux t6237 (
    .I(seg_16_14_sp4_h_r_8_66015),
    .O(seg_16_14_local_g0_0_65911)
  );
  LocalMux t6238 (
    .I(seg_16_14_sp4_h_r_12_62175),
    .O(seg_16_14_local_g1_4_65923)
  );
  LocalMux t6239 (
    .I(seg_16_14_sp4_h_r_14_62179),
    .O(seg_16_14_local_g1_6_65925)
  );
  CascadeMux t624 (
    .I(net_46553),
    .O(net_46553_cascademuxed)
  );
  LocalMux t6240 (
    .I(seg_16_14_sp4_h_r_16_62181),
    .O(seg_16_14_local_g1_0_65919)
  );
  LocalMux t6241 (
    .I(seg_18_10_sp4_h_r_40_61689),
    .O(seg_18_10_local_g2_0_73097)
  );
  Span4Mux_h1 t6242 (
    .I(seg_19_10_sp4_v_t_46_73320),
    .O(seg_18_10_sp4_h_r_40_61689)
  );
  LocalMux t6243 (
    .I(seg_18_10_sp4_v_b_17_69115),
    .O(seg_18_10_local_g0_1_73082)
  );
  Span4Mux_v1 t6244 (
    .I(seg_18_11_sp4_v_t_36_69602),
    .O(seg_18_10_sp4_v_b_17_69115)
  );
  LocalMux t6245 (
    .I(seg_17_16_neigh_op_bnr_1_69825),
    .O(seg_17_16_local_g1_1_69997)
  );
  LocalMux t6246 (
    .I(seg_17_16_neigh_op_bnr_2_69826),
    .O(seg_17_16_local_g0_2_69990)
  );
  LocalMux t6247 (
    .I(seg_17_16_neigh_op_bnr_3_69827),
    .O(seg_17_16_local_g0_3_69991)
  );
  LocalMux t6248 (
    .I(seg_17_16_neigh_op_bnr_4_69828),
    .O(seg_17_16_local_g1_4_70000)
  );
  LocalMux t6249 (
    .I(seg_17_16_neigh_op_bnr_5_69829),
    .O(seg_17_16_local_g1_5_70001)
  );
  CascadeMux t625 (
    .I(net_46571),
    .O(net_46571_cascademuxed)
  );
  LocalMux t6250 (
    .I(seg_17_16_neigh_op_bnr_6_69830),
    .O(seg_17_16_local_g1_6_70002)
  );
  LocalMux t6251 (
    .I(seg_17_16_neigh_op_bnr_7_69831),
    .O(seg_17_16_local_g1_7_70003)
  );
  LocalMux t6252 (
    .I(seg_17_17_neigh_op_bnr_0_69947),
    .O(seg_17_17_local_g0_0_70111)
  );
  LocalMux t6253 (
    .I(seg_18_16_lutff_1_out_69948),
    .O(seg_18_16_local_g3_1_73844)
  );
  LocalMux t6254 (
    .I(seg_17_15_neigh_op_tnr_2_69949),
    .O(seg_17_15_local_g2_2_69883)
  );
  LocalMux t6255 (
    .I(seg_18_15_neigh_op_top_2_69949),
    .O(seg_18_15_local_g1_2_73706)
  );
  LocalMux t6256 (
    .I(seg_17_16_neigh_op_rgt_4_69951),
    .O(seg_17_16_local_g3_4_70016)
  );
  LocalMux t6257 (
    .I(seg_17_17_neigh_op_bnr_4_69951),
    .O(seg_17_17_local_g0_4_70115)
  );
  LocalMux t6258 (
    .I(seg_17_15_neigh_op_tnr_5_69952),
    .O(seg_17_15_local_g2_5_69886)
  );
  LocalMux t6259 (
    .I(seg_18_15_neigh_op_top_5_69952),
    .O(seg_18_15_local_g1_5_73709)
  );
  CascadeMux t626 (
    .I(net_46577),
    .O(net_46577_cascademuxed)
  );
  LocalMux t6260 (
    .I(seg_16_15_sp4_v_b_14_62065),
    .O(seg_16_15_local_g0_6_66040)
  );
  Span4Mux_v1 t6261 (
    .I(seg_16_16_sp4_h_r_10_66253),
    .O(seg_16_15_sp4_v_b_14_62065)
  );
  LocalMux t6262 (
    .I(seg_18_13_sp4_v_b_47_69736),
    .O(seg_18_13_local_g3_7_73481)
  );
  LocalMux t6263 (
    .I(seg_17_12_sp4_r_v_b_5_69237),
    .O(seg_17_12_local_g1_5_69509)
  );
  Span4Mux_v1 t6264 (
    .I(seg_18_12_sp4_v_t_39_69728),
    .O(seg_17_12_sp4_r_v_b_5_69237)
  );
  LocalMux t6265 (
    .I(seg_16_14_sp4_h_r_30_58352),
    .O(seg_16_14_local_g2_6_65933)
  );
  Span4Mux_h2 t6266 (
    .I(seg_18_14_sp4_v_t_43_69978),
    .O(seg_16_14_sp4_h_r_30_58352)
  );
  LocalMux t6267 (
    .I(seg_18_15_sp4_v_b_43_69978),
    .O(seg_18_15_local_g3_3_73723)
  );
  LocalMux t6268 (
    .I(seg_18_13_sp4_v_b_41_69730),
    .O(seg_18_13_local_g2_1_73467)
  );
  LocalMux t6269 (
    .I(seg_17_16_neigh_op_tnr_4_70074),
    .O(seg_17_16_local_g2_4_70008)
  );
  CascadeMux t627 (
    .I(net_46682),
    .O(net_46682_cascademuxed)
  );
  LocalMux t6270 (
    .I(seg_17_17_neigh_op_rgt_4_70074),
    .O(seg_17_17_local_g2_4_70131)
  );
  GlobalMux t6271 (
    .I(seg_13_0_local_g1_4_52735_i3),
    .O(seg_1_1_glb_netwk_0_5)
  );
  gio2CtrlBuf t6272 (
    .I(seg_13_0_local_g1_4_52735_i2),
    .O(seg_13_0_local_g1_4_52735_i3)
  );
  ICE_GB t6273 (
    .GLOBALBUFFEROUTPUT(seg_13_0_local_g1_4_52735_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_13_0_local_g1_4_52735_i1)
  );
  IoInMux t6274 (
    .I(seg_13_0_local_g1_4_52735),
    .O(seg_13_0_local_g1_4_52735_i1)
  );
  LocalMux t6275 (
    .I(seg_13_0_span4_horz_r_4_48940),
    .O(seg_13_0_local_g1_4_52735)
  );
  IoSpan4Mux t6276 (
    .I(seg_16_0_span4_horz_r_0_64262),
    .O(seg_13_0_span4_horz_r_4_48940)
  );
  LocalMux t6277 (
    .I(seg_3_2_sp4_h_r_7_15368),
    .O(seg_3_2_local_g1_7_15280)
  );
  Span4Mux_h4 t6278 (
    .I(seg_7_2_sp4_h_r_4_30058),
    .O(seg_3_2_sp4_h_r_7_15368)
  );
  Span4Mux_h4 t6279 (
    .I(seg_11_2_sp4_h_r_4_45382),
    .O(seg_7_2_sp4_h_r_4_30058)
  );
  CascadeMux t628 (
    .I(net_46694),
    .O(net_46694_cascademuxed)
  );
  Span4Mux_h4 t6280 (
    .I(seg_15_2_sp4_h_r_1_60699),
    .O(seg_11_2_sp4_h_r_4_45382)
  );
  Span4Mux_h4 t6281 (
    .I(seg_19_2_sp4_v_b_1_72048),
    .O(seg_15_2_sp4_h_r_1_60699)
  );
  LocalMux t6282 (
    .I(seg_4_2_sp4_h_r_13_15359),
    .O(seg_4_2_local_g1_5_19109)
  );
  Span4Mux_h3 t6283 (
    .I(seg_7_2_sp4_h_r_4_30058),
    .O(seg_4_2_sp4_h_r_13_15359)
  );
  LocalMux t6284 (
    .I(seg_20_2_lutff_2_out_75801),
    .O(seg_20_2_local_g0_2_79130)
  );
  LocalMux t6285 (
    .I(seg_20_2_lutff_7_out_75806),
    .O(seg_20_2_local_g1_7_79143)
  );
  LocalMux t6286 (
    .I(seg_18_2_sp4_h_r_12_68361),
    .O(seg_18_2_local_g1_4_72109)
  );
  LocalMux t6287 (
    .I(seg_18_2_sp4_h_r_22_68363),
    .O(seg_18_2_local_g0_6_72103)
  );
  LocalMux t6288 (
    .I(seg_20_3_lutff_0_out_75937),
    .O(seg_20_3_local_g1_0_79259)
  );
  LocalMux t6289 (
    .I(seg_20_3_lutff_1_out_75938),
    .O(seg_20_3_local_g2_1_79268)
  );
  CascadeMux t629 (
    .I(net_46817),
    .O(net_46817_cascademuxed)
  );
  LocalMux t6290 (
    .I(seg_18_3_sp4_h_r_4_72320),
    .O(seg_18_3_local_g0_4_72224)
  );
  LocalMux t6291 (
    .I(seg_17_3_sp4_h_r_3_68488),
    .O(seg_17_3_local_g1_3_68400)
  );
  LocalMux t6292 (
    .I(seg_18_3_sp4_h_r_18_68492),
    .O(seg_18_3_local_g0_2_72222)
  );
  LocalMux t6293 (
    .I(seg_17_3_sp4_h_r_11_68486),
    .O(seg_17_3_local_g0_3_68392)
  );
  LocalMux t6294 (
    .I(seg_23_0_span4_vert_42_86774),
    .O(seg_23_0_local_g1_2_90410)
  );
  Span4Mux_v4 t6295 (
    .I(seg_23_4_sp4_h_l_42_76192),
    .O(seg_23_0_span4_vert_42_86774)
  );
  LocalMux t6296 (
    .I(seg_18_9_sp4_h_r_15_69225),
    .O(seg_18_9_local_g1_7_72973)
  );
  Span4Mux_h3 t6297 (
    .I(seg_21_9_sp4_v_b_9_79734),
    .O(seg_18_9_sp4_h_r_15_69225)
  );
  Span4Mux_v4 t6298 (
    .I(seg_21_5_sp4_v_b_6_79241),
    .O(seg_21_9_sp4_v_b_9_79734)
  );
  LocalMux t6299 (
    .I(seg_16_5_sp4_h_r_16_61074),
    .O(seg_16_5_local_g1_0_64812)
  );
  CascadeMux t63 (
    .I(net_11481),
    .O(net_11481_cascademuxed)
  );
  CascadeMux t630 (
    .I(net_46928),
    .O(net_46928_cascademuxed)
  );
  Span4Mux_h3 t6300 (
    .I(seg_19_5_sp4_h_r_5_76292),
    .O(seg_16_5_sp4_h_r_16_61074)
  );
  LocalMux t6301 (
    .I(seg_17_5_sp4_h_r_15_64902),
    .O(seg_17_5_local_g0_7_68642)
  );
  Span4Mux_h3 t6302 (
    .I(seg_20_5_sp4_h_r_2_79595),
    .O(seg_17_5_sp4_h_r_15_64902)
  );
  LocalMux t6303 (
    .I(seg_18_5_sp4_h_r_4_72566),
    .O(seg_18_5_local_g0_4_72470)
  );
  LocalMux t6304 (
    .I(seg_17_5_sp4_h_r_1_68730),
    .O(seg_17_5_local_g1_1_68644)
  );
  LocalMux t6305 (
    .I(seg_17_5_sp4_h_r_3_68734),
    .O(seg_17_5_local_g1_3_68646)
  );
  LocalMux t6306 (
    .I(seg_16_5_sp4_r_v_b_5_64545),
    .O(seg_16_5_local_g1_5_64817)
  );
  Span4Mux_v1 t6307 (
    .I(seg_17_5_sp4_h_r_5_68736),
    .O(seg_16_5_sp4_r_v_b_5_64545)
  );
  LocalMux t6308 (
    .I(seg_17_4_sp4_v_b_18_64547),
    .O(seg_17_4_local_g1_2_68522)
  );
  Span4Mux_v1 t6309 (
    .I(seg_17_5_sp4_h_r_7_68738),
    .O(seg_17_4_sp4_v_b_18_64547)
  );
  CascadeMux t631 (
    .I(net_46958),
    .O(net_46958_cascademuxed)
  );
  LocalMux t6310 (
    .I(seg_17_5_sp4_h_r_11_68732),
    .O(seg_17_5_local_g0_3_68638)
  );
  LocalMux t6311 (
    .I(seg_18_6_sp4_h_r_8_72693),
    .O(seg_18_6_local_g1_0_72597)
  );
  LocalMux t6312 (
    .I(seg_17_6_sp4_h_r_5_68859),
    .O(seg_17_6_local_g1_5_68771)
  );
  LocalMux t6313 (
    .I(seg_15_7_sp4_r_v_b_15_61082),
    .O(seg_15_7_local_g2_7_61242)
  );
  Span4Mux_v1 t6314 (
    .I(seg_16_8_sp4_h_r_2_65271),
    .O(seg_15_7_sp4_r_v_b_15_61082)
  );
  Span4Mux_h4 t6315 (
    .I(seg_20_8_sp4_v_b_2_76300),
    .O(seg_16_8_sp4_h_r_2_65271)
  );
  LocalMux t6316 (
    .I(seg_15_7_sp4_h_r_27_53658),
    .O(seg_15_7_local_g3_3_61246)
  );
  Span4Mux_h2 t6317 (
    .I(seg_17_7_sp4_h_r_7_68984),
    .O(seg_15_7_sp4_h_r_27_53658)
  );
  LocalMux t6318 (
    .I(seg_16_8_sp4_h_r_20_61447),
    .O(seg_16_8_local_g1_4_65185)
  );
  Span4Mux_h3 t6319 (
    .I(seg_19_8_sp4_h_r_1_76592),
    .O(seg_16_8_sp4_h_r_20_61447)
  );
  CascadeMux t632 (
    .I(net_47039),
    .O(net_47039_cascademuxed)
  );
  LocalMux t6320 (
    .I(seg_16_6_sp4_h_r_10_65023),
    .O(seg_16_6_local_g0_2_64929)
  );
  Span4Mux_h4 t6321 (
    .I(seg_20_6_sp4_v_t_41_76506),
    .O(seg_16_6_sp4_h_r_10_65023)
  );
  LocalMux t6322 (
    .I(seg_20_10_neigh_op_bot_7_76556),
    .O(seg_20_10_local_g0_7_80119)
  );
  LocalMux t6323 (
    .I(seg_16_9_sp4_r_v_b_0_65034),
    .O(seg_16_9_local_g1_0_65304)
  );
  Span4Mux_v1 t6324 (
    .I(seg_17_9_sp4_h_r_7_69230),
    .O(seg_16_9_sp4_r_v_b_0_65034)
  );
  LocalMux t6325 (
    .I(seg_16_9_sp4_h_r_11_65393),
    .O(seg_16_9_local_g1_3_65307)
  );
  Span4Mux_h4 t6326 (
    .I(seg_20_9_sp4_h_r_8_80093),
    .O(seg_16_9_sp4_h_r_11_65393)
  );
  LocalMux t6327 (
    .I(seg_12_10_sp4_h_r_11_50194),
    .O(seg_12_10_local_g1_3_50108)
  );
  Span4Mux_h4 t6328 (
    .I(seg_16_10_sp4_h_r_11_65516),
    .O(seg_12_10_sp4_h_r_11_50194)
  );
  Span4Mux_h4 t6329 (
    .I(seg_20_10_sp4_v_b_11_76511),
    .O(seg_16_10_sp4_h_r_11_65516)
  );
  CascadeMux t633 (
    .I(net_47045),
    .O(net_47045_cascademuxed)
  );
  LocalMux t6330 (
    .I(seg_21_10_neigh_op_lft_0_76651),
    .O(seg_21_10_local_g0_0_83943)
  );
  LocalMux t6331 (
    .I(seg_20_11_neigh_op_bot_1_76652),
    .O(seg_20_11_local_g1_1_80244)
  );
  LocalMux t6332 (
    .I(seg_21_10_neigh_op_lft_5_76656),
    .O(seg_21_10_local_g1_5_83956)
  );
  LocalMux t6333 (
    .I(seg_18_9_sp4_v_b_13_68988),
    .O(seg_18_9_local_g1_5_72971)
  );
  Span4Mux_v1 t6334 (
    .I(seg_18_10_sp4_h_r_0_73175),
    .O(seg_18_9_sp4_v_b_13_68988)
  );
  LocalMux t6335 (
    .I(seg_22_0_span4_vert_22_82921),
    .O(seg_22_0_local_g1_6_86583)
  );
  Span4Mux_v2 t6336 (
    .I(seg_22_2_sp4_v_t_46_83198),
    .O(seg_22_0_span4_vert_22_82921)
  );
  Span4Mux_v4 t6337 (
    .I(seg_22_6_sp4_v_t_45_83689),
    .O(seg_22_2_sp4_v_t_46_83198)
  );
  Span4Mux_v4 t6338 (
    .I(seg_22_10_sp4_h_l_39_73179),
    .O(seg_22_6_sp4_v_t_45_83689)
  );
  LocalMux t6339 (
    .I(seg_20_10_neigh_op_top_6_76759),
    .O(seg_20_10_local_g1_6_80126)
  );
  CascadeMux t634 (
    .I(net_47057),
    .O(net_47057_cascademuxed)
  );
  LocalMux t6340 (
    .I(seg_18_10_sp4_v_b_22_69120),
    .O(seg_18_10_local_g1_6_73095)
  );
  Span4Mux_v1 t6341 (
    .I(seg_18_11_sp4_h_r_6_73306),
    .O(seg_18_10_sp4_v_b_22_69120)
  );
  LocalMux t6342 (
    .I(seg_13_8_sp4_h_r_18_49954),
    .O(seg_13_8_local_g1_2_53692)
  );
  Span4Mux_h3 t6343 (
    .I(seg_16_8_sp4_h_r_4_65273),
    .O(seg_13_8_sp4_h_r_18_49954)
  );
  Span4Mux_h4 t6344 (
    .I(seg_20_8_sp4_v_t_41_76710),
    .O(seg_16_8_sp4_h_r_4_65273)
  );
  LocalMux t6345 (
    .I(seg_13_14_sp4_h_r_3_54519),
    .O(seg_13_14_local_g1_3_54431)
  );
  Span4Mux_h4 t6346 (
    .I(seg_17_14_sp4_h_r_3_69841),
    .O(seg_13_14_sp4_h_r_3_54519)
  );
  LocalMux t6347 (
    .I(seg_20_3_neigh_op_rgt_3_79213),
    .O(seg_20_3_local_g3_3_79278)
  );
  LocalMux t6348 (
    .I(seg_18_3_sp4_h_r_21_68493),
    .O(seg_18_3_local_g1_5_72233)
  );
  Span4Mux_h3 t6349 (
    .I(seg_21_3_sp4_h_r_0_83176),
    .O(seg_18_3_sp4_h_r_21_68493)
  );
  CascadeMux t635 (
    .I(net_47063),
    .O(net_47063_cascademuxed)
  );
  LocalMux t6350 (
    .I(seg_18_3_sp4_h_r_1_72315),
    .O(seg_18_3_local_g1_1_72229)
  );
  LocalMux t6351 (
    .I(seg_18_3_sp4_h_r_11_72317),
    .O(seg_18_3_local_g0_3_72223)
  );
  LocalMux t6352 (
    .I(seg_17_4_sp4_h_r_21_64785),
    .O(seg_17_4_local_g1_5_68525)
  );
  Span4Mux_h3 t6353 (
    .I(seg_20_4_sp4_h_r_5_79475),
    .O(seg_17_4_sp4_h_r_21_64785)
  );
  LocalMux t6354 (
    .I(seg_17_4_sp4_h_r_23_64777),
    .O(seg_17_4_local_g1_7_68527)
  );
  Span4Mux_h3 t6355 (
    .I(seg_20_4_sp4_h_r_7_79477),
    .O(seg_17_4_sp4_h_r_23_64777)
  );
  LocalMux t6356 (
    .I(seg_18_4_sp4_h_r_1_72438),
    .O(seg_18_4_local_g1_1_72352)
  );
  LocalMux t6357 (
    .I(seg_17_4_sp4_r_v_b_0_68244),
    .O(seg_17_4_local_g1_0_68520)
  );
  Span4Mux_v1 t6358 (
    .I(seg_18_4_sp4_h_r_7_72446),
    .O(seg_17_4_sp4_r_v_b_0_68244)
  );
  LocalMux t6359 (
    .I(seg_18_4_sp4_h_r_11_72440),
    .O(seg_18_4_local_g1_3_72354)
  );
  LocalMux t6360 (
    .I(seg_18_5_sp4_h_r_1_72561),
    .O(seg_18_5_local_g1_1_72475)
  );
  LocalMux t6361 (
    .I(seg_17_5_sp4_r_v_b_10_68383),
    .O(seg_17_5_local_g2_2_68653)
  );
  Span4Mux_v1 t6362 (
    .I(seg_18_5_sp4_h_r_5_72567),
    .O(seg_17_5_sp4_r_v_b_10_68383)
  );
  LocalMux t6363 (
    .I(seg_17_4_sp4_r_v_b_15_68375),
    .O(seg_17_4_local_g2_7_68535)
  );
  Span4Mux_v1 t6364 (
    .I(seg_18_5_sp4_h_r_9_72571),
    .O(seg_17_4_sp4_r_v_b_15_68375)
  );
  LocalMux t6365 (
    .I(seg_21_6_lutff_6_out_79585),
    .O(seg_21_6_local_g3_6_83481)
  );
  LocalMux t6366 (
    .I(seg_17_6_sp4_h_r_22_65024),
    .O(seg_17_6_local_g0_6_68764)
  );
  Span4Mux_h3 t6367 (
    .I(seg_20_6_sp4_h_r_3_79719),
    .O(seg_17_6_sp4_h_r_22_65024)
  );
  LocalMux t6368 (
    .I(seg_18_5_sp4_v_b_16_68499),
    .O(seg_18_5_local_g1_0_72474)
  );
  Span4Mux_v1 t6369 (
    .I(seg_18_6_sp4_h_r_5_72690),
    .O(seg_18_5_sp4_v_b_16_68499)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t637 (
    .carryinitin(),
    .carryinitout(t636)
  );
  LocalMux t6370 (
    .I(seg_18_6_sp4_h_r_7_72692),
    .O(seg_18_6_local_g1_7_72604)
  );
  LocalMux t6371 (
    .I(seg_21_8_neigh_op_bot_1_79703),
    .O(seg_21_8_local_g1_1_83706)
  );
  LocalMux t6372 (
    .I(seg_21_8_neigh_op_bot_2_79704),
    .O(seg_21_8_local_g0_2_83699)
  );
  LocalMux t6373 (
    .I(seg_18_6_sp4_v_b_21_68627),
    .O(seg_18_6_local_g0_5_72594)
  );
  Span4Mux_v1 t6374 (
    .I(seg_18_7_sp4_h_r_3_72811),
    .O(seg_18_6_sp4_v_b_21_68627)
  );
  LocalMux t6375 (
    .I(seg_17_6_sp4_r_v_b_17_68623),
    .O(seg_17_6_local_g3_1_68783)
  );
  Span4Mux_v1 t6376 (
    .I(seg_18_7_sp4_h_r_11_72809),
    .O(seg_17_6_sp4_r_v_b_17_68623)
  );
  LocalMux t6377 (
    .I(seg_20_9_neigh_op_bnr_1_79826),
    .O(seg_20_9_local_g1_1_79998)
  );
  LocalMux t6378 (
    .I(seg_20_9_neigh_op_bnr_7_79832),
    .O(seg_20_9_local_g1_7_80004)
  );
  LocalMux t6379 (
    .I(seg_16_8_sp12_h_r_3_61432),
    .O(seg_16_8_local_g0_3_65176)
  );
  LocalMux t6380 (
    .I(seg_16_8_sp12_h_r_5_57603),
    .O(seg_16_8_local_g1_5_65186)
  );
  LocalMux t6381 (
    .I(seg_18_8_sp4_h_r_5_72936),
    .O(seg_18_8_local_g1_5_72848)
  );
  LocalMux t6382 (
    .I(seg_18_8_sp4_h_r_9_72940),
    .O(seg_18_8_local_g0_1_72836)
  );
  LocalMux t6383 (
    .I(seg_16_9_sp4_r_v_b_15_65159),
    .O(seg_16_9_local_g2_7_65319)
  );
  Span4Mux_v1 t6384 (
    .I(seg_17_10_sp4_h_r_2_69348),
    .O(seg_16_9_sp4_r_v_b_15_65159)
  );
  Span4Mux_h4 t6385 (
    .I(seg_21_10_sp4_v_b_2_79852),
    .O(seg_17_10_sp4_h_r_2_69348)
  );
  LocalMux t6386 (
    .I(seg_21_10_neigh_op_bot_0_79948),
    .O(seg_21_10_local_g1_0_83951)
  );
  LocalMux t6387 (
    .I(seg_20_8_neigh_op_tnr_3_79951),
    .O(seg_20_8_local_g3_3_79893)
  );
  LocalMux t6388 (
    .I(seg_21_9_lutff_4_out_79952),
    .O(seg_21_9_local_g1_4_83832)
  );
  LocalMux t6389 (
    .I(seg_21_8_neigh_op_top_6_79954),
    .O(seg_21_8_local_g1_6_83711)
  );
  CascadeMux t639 (
    .I(net_47162),
    .O(net_47162_cascademuxed)
  );
  LocalMux t6390 (
    .I(seg_21_9_lutff_6_out_79954),
    .O(seg_21_9_local_g3_6_83850)
  );
  LocalMux t6391 (
    .I(seg_20_9_neigh_op_rgt_7_79955),
    .O(seg_20_9_local_g3_7_80020)
  );
  LocalMux t6392 (
    .I(seg_17_9_sp4_h_r_20_65401),
    .O(seg_17_9_local_g0_4_69131)
  );
  Span4Mux_h3 t6393 (
    .I(seg_20_9_sp4_h_r_9_80094),
    .O(seg_17_9_sp4_h_r_20_65401)
  );
  LocalMux t6394 (
    .I(seg_17_10_sp4_h_r_0_69344),
    .O(seg_17_10_local_g1_0_69258)
  );
  Span4Mux_h4 t6395 (
    .I(seg_21_10_sp4_v_b_7_79855),
    .O(seg_17_10_sp4_h_r_0_69344)
  );
  LocalMux t6396 (
    .I(seg_21_9_neigh_op_top_2_80073),
    .O(seg_21_9_local_g1_2_83830)
  );
  LocalMux t6397 (
    .I(seg_21_9_neigh_op_top_3_80074),
    .O(seg_21_9_local_g1_3_83831)
  );
  LocalMux t6398 (
    .I(seg_18_10_sp4_h_r_21_69354),
    .O(seg_18_10_local_g0_5_73086)
  );
  Span4Mux_h3 t6399 (
    .I(seg_21_10_sp4_h_r_0_84037),
    .O(seg_18_10_sp4_h_r_21_69354)
  );
  CascadeMux t64 (
    .I(net_11487),
    .O(net_11487_cascademuxed)
  );
  CascadeMux t640 (
    .I(net_47192),
    .O(net_47192_cascademuxed)
  );
  LocalMux t6400 (
    .I(seg_18_10_sp4_h_r_16_69351),
    .O(seg_18_10_local_g0_0_73081)
  );
  Span4Mux_h3 t6401 (
    .I(seg_21_10_sp4_h_r_2_84041),
    .O(seg_18_10_sp4_h_r_16_69351)
  );
  LocalMux t6402 (
    .I(seg_18_11_sp4_v_b_40_69483),
    .O(seg_18_11_local_g3_0_73228)
  );
  Span4Mux_v1 t6403 (
    .I(seg_18_10_sp4_h_r_5_73182),
    .O(seg_18_11_sp4_v_b_40_69483)
  );
  LocalMux t6404 (
    .I(seg_21_3_neigh_op_rgt_0_83041),
    .O(seg_21_3_local_g3_0_83106)
  );
  LocalMux t6405 (
    .I(seg_21_3_neigh_op_rgt_2_83043),
    .O(seg_21_3_local_g2_2_83100)
  );
  LocalMux t6406 (
    .I(seg_18_3_sp4_h_r_8_72324),
    .O(seg_18_3_local_g1_0_72228)
  );
  Span4Mux_h4 t6407 (
    .I(seg_22_3_sp4_h_r_8_87017),
    .O(seg_18_3_sp4_h_r_8_72324)
  );
  LocalMux t6408 (
    .I(seg_21_3_neigh_op_tnr_6_83170),
    .O(seg_21_3_local_g3_6_83112)
  );
  LocalMux t6409 (
    .I(seg_21_4_neigh_op_rgt_7_83171),
    .O(seg_21_4_local_g2_7_83228)
  );
  CascadeMux t641 (
    .I(net_47198),
    .O(net_47198_cascademuxed)
  );
  LocalMux t6410 (
    .I(seg_17_4_sp12_h_r_3_64771),
    .O(seg_17_4_local_g1_3_68523)
  );
  LocalMux t6411 (
    .I(seg_21_5_neigh_op_rgt_4_83291),
    .O(seg_21_5_local_g3_4_83356)
  );
  LocalMux t6412 (
    .I(seg_21_4_neigh_op_tnr_6_83293),
    .O(seg_21_4_local_g2_6_83227)
  );
  LocalMux t6413 (
    .I(seg_18_5_sp4_h_r_19_68737),
    .O(seg_18_5_local_g1_3_72477)
  );
  Span4Mux_h3 t6414 (
    .I(seg_21_5_sp4_h_r_3_83427),
    .O(seg_18_5_sp4_h_r_19_68737)
  );
  LocalMux t6415 (
    .I(seg_20_5_sp4_h_r_8_79601),
    .O(seg_20_5_local_g1_0_79505)
  );
  LocalMux t6416 (
    .I(seg_18_5_sp4_r_v_b_8_72212),
    .O(seg_18_5_local_g2_0_72482)
  );
  Span4Mux_v1 t6417 (
    .I(seg_19_5_sp4_h_r_3_76290),
    .O(seg_18_5_sp4_r_v_b_8_72212)
  );
  LocalMux t6418 (
    .I(seg_21_6_neigh_op_rgt_4_83414),
    .O(seg_21_6_local_g3_4_83479)
  );
  LocalMux t6419 (
    .I(seg_18_6_sp4_h_r_17_68858),
    .O(seg_18_6_local_g1_1_72598)
  );
  CascadeMux t642 (
    .I(net_47291),
    .O(net_47291_cascademuxed)
  );
  Span4Mux_h3 t6420 (
    .I(seg_21_6_sp4_h_r_1_83546),
    .O(seg_18_6_sp4_h_r_17_68858)
  );
  LocalMux t6421 (
    .I(seg_21_8_neigh_op_bnr_2_83535),
    .O(seg_21_8_local_g1_2_83707)
  );
  LocalMux t6422 (
    .I(seg_21_8_neigh_op_bnr_4_83537),
    .O(seg_21_8_local_g0_4_83701)
  );
  LocalMux t6423 (
    .I(seg_21_8_neigh_op_bnr_5_83538),
    .O(seg_21_8_local_g1_5_83710)
  );
  LocalMux t6424 (
    .I(seg_21_8_neigh_op_bnr_7_83540),
    .O(seg_21_8_local_g0_7_83704)
  );
  LocalMux t6425 (
    .I(seg_21_8_neigh_op_rgt_0_83656),
    .O(seg_21_8_local_g3_0_83721)
  );
  LocalMux t6426 (
    .I(seg_21_7_neigh_op_tnr_2_83658),
    .O(seg_21_7_local_g3_2_83600)
  );
  LocalMux t6427 (
    .I(seg_21_8_neigh_op_rgt_3_83659),
    .O(seg_21_8_local_g2_3_83716)
  );
  LocalMux t6428 (
    .I(seg_21_8_neigh_op_rgt_4_83660),
    .O(seg_21_8_local_g2_4_83717)
  );
  LocalMux t6429 (
    .I(seg_21_8_neigh_op_rgt_5_83661),
    .O(seg_21_8_local_g3_5_83726)
  );
  CascadeMux t643 (
    .I(net_47297),
    .O(net_47297_cascademuxed)
  );
  LocalMux t6430 (
    .I(seg_21_9_neigh_op_bnr_5_83661),
    .O(seg_21_9_local_g0_5_83825)
  );
  LocalMux t6431 (
    .I(seg_21_8_neigh_op_rgt_6_83662),
    .O(seg_21_8_local_g2_6_83719)
  );
  LocalMux t6432 (
    .I(seg_21_9_neigh_op_rgt_0_83779),
    .O(seg_21_9_local_g2_0_83836)
  );
  LocalMux t6433 (
    .I(seg_21_9_neigh_op_rgt_3_83782),
    .O(seg_21_9_local_g3_3_83847)
  );
  LocalMux t6434 (
    .I(seg_21_8_neigh_op_tnr_4_83783),
    .O(seg_21_8_local_g3_4_83725)
  );
  LocalMux t6435 (
    .I(seg_21_8_neigh_op_tnr_6_83785),
    .O(seg_21_8_local_g3_6_83727)
  );
  LocalMux t6436 (
    .I(seg_21_8_neigh_op_tnr_7_83786),
    .O(seg_21_8_local_g2_7_83720)
  );
  LocalMux t6437 (
    .I(seg_17_10_sp4_h_r_21_65523),
    .O(seg_17_10_local_g1_5_69263)
  );
  Span4Mux_h3 t6438 (
    .I(seg_20_10_sp4_h_r_8_80216),
    .O(seg_17_10_sp4_h_r_21_65523)
  );
  LocalMux t6439 (
    .I(seg_3_1_sp4_h_r_4_15206),
    .O(seg_3_1_local_g0_4_15106)
  );
  CascadeMux t644 (
    .I(net_47315),
    .O(net_47315_cascademuxed)
  );
  Span4Mux_h4 t6440 (
    .I(seg_7_1_sp4_h_r_8_29903),
    .O(seg_3_1_sp4_h_r_4_15206)
  );
  Span4Mux_h4 t6441 (
    .I(seg_11_1_sp4_h_r_8_45227),
    .O(seg_7_1_sp4_h_r_8_29903)
  );
  Span4Mux_h4 t6442 (
    .I(seg_15_1_sp4_h_r_5_60546),
    .O(seg_11_1_sp4_h_r_8_45227)
  );
  Span4Mux_h4 t6443 (
    .I(seg_19_1_sp4_h_r_5_75848),
    .O(seg_15_1_sp4_h_r_5_60546)
  );
  Span4Mux_h4 t6444 (
    .I(seg_23_1_sp4_v_b_0_86737),
    .O(seg_19_1_sp4_h_r_5_75848)
  );
  LocalMux t6445 (
    .I(seg_4_2_sp4_h_r_14_15364),
    .O(seg_4_2_local_g1_6_19110)
  );
  Span4Mux_h3 t6446 (
    .I(seg_7_2_sp4_h_r_7_30061),
    .O(seg_4_2_sp4_h_r_14_15364)
  );
  Span4Mux_h4 t6447 (
    .I(seg_11_2_sp4_h_r_11_45379),
    .O(seg_7_2_sp4_h_r_7_30061)
  );
  Span4Mux_h4 t6448 (
    .I(seg_15_2_sp4_h_r_8_60708),
    .O(seg_11_2_sp4_h_r_11_45379)
  );
  Span4Mux_h4 t6449 (
    .I(seg_19_2_sp4_h_r_5_75986),
    .O(seg_15_2_sp4_h_r_8_60708)
  );
  CascadeMux t645 (
    .I(net_47327),
    .O(net_47327_cascademuxed)
  );
  Span4Mux_h4 t6450 (
    .I(seg_23_2_sp4_v_b_5_86745),
    .O(seg_19_2_sp4_h_r_5_75986)
  );
  LocalMux t6451 (
    .I(seg_22_5_neigh_op_rgt_0_87118),
    .O(seg_22_5_local_g3_0_87183)
  );
  LocalMux t6452 (
    .I(seg_22_5_neigh_op_rgt_1_87119),
    .O(seg_22_5_local_g2_1_87176)
  );
  LocalMux t6453 (
    .I(seg_22_4_neigh_op_tnr_7_87125),
    .O(seg_22_4_local_g2_7_87059)
  );
  LocalMux t6454 (
    .I(seg_17_5_sp4_h_r_16_64905),
    .O(seg_17_5_local_g1_0_68643)
  );
  Span4Mux_h3 t6455 (
    .I(seg_20_5_sp4_h_r_5_79598),
    .O(seg_17_5_sp4_h_r_16_64905)
  );
  LocalMux t6456 (
    .I(seg_18_3_sp4_r_v_b_7_72069),
    .O(seg_18_3_local_g1_7_72235)
  );
  Span4Mux_v1 t6457 (
    .I(seg_19_3_sp4_h_r_2_76085),
    .O(seg_18_3_sp4_r_v_b_7_72069)
  );
  Span4Mux_h4 t6458 (
    .I(seg_23_3_sp4_v_t_39_87145),
    .O(seg_19_3_sp4_h_r_2_76085)
  );
  LocalMux t6459 (
    .I(seg_23_5_neigh_op_top_1_87242),
    .O(seg_23_5_local_g0_1_90991)
  );
  CascadeMux t646 (
    .I(net_48985),
    .O(net_48985_cascademuxed)
  );
  LocalMux t6460 (
    .I(seg_22_5_neigh_op_tnr_3_87244),
    .O(seg_22_5_local_g2_3_87178)
  );
  LocalMux t6461 (
    .I(seg_22_6_neigh_op_rgt_7_87248),
    .O(seg_22_6_local_g2_7_87305)
  );
  LocalMux t6462 (
    .I(seg_21_8_sp4_h_r_6_83799),
    .O(seg_21_8_local_g0_6_83703)
  );
  LocalMux t6463 (
    .I(seg_21_9_sp4_h_r_14_80088),
    .O(seg_21_9_local_g1_6_83834)
  );
  LocalMux t6464 (
    .I(seg_22_7_sp4_r_v_b_24_87389),
    .O(seg_22_7_local_g1_0_87413)
  );
  Span4Mux_v2 t6465 (
    .I(seg_23_5_sp4_h_r_0_91084),
    .O(seg_22_7_sp4_r_v_b_24_87389)
  );
  LocalMux t6466 (
    .I(seg_22_8_sp4_r_v_b_21_87397),
    .O(seg_22_8_local_g3_5_87557)
  );
  Span4Mux_v3 t6467 (
    .I(seg_23_5_sp4_h_r_8_91094),
    .O(seg_22_8_sp4_r_v_b_21_87397)
  );
  LocalMux t6468 (
    .I(seg_22_7_sp4_v_b_31_83563),
    .O(seg_22_7_local_g2_7_87428)
  );
  Span4Mux_v2 t6469 (
    .I(seg_22_5_sp4_h_r_1_87254),
    .O(seg_22_7_sp4_v_b_31_83563)
  );
  CascadeMux t647 (
    .I(net_48997),
    .O(net_48997_cascademuxed)
  );
  LocalMux t6470 (
    .I(seg_21_7_sp4_r_v_b_33_83565),
    .O(seg_21_7_local_g0_2_83576)
  );
  Span4Mux_v2 t6471 (
    .I(seg_22_5_sp4_h_r_3_87258),
    .O(seg_21_7_sp4_r_v_b_33_83565)
  );
  LocalMux t6472 (
    .I(seg_22_7_sp4_v_b_25_83557),
    .O(seg_22_7_local_g3_1_87430)
  );
  Span4Mux_v2 t6473 (
    .I(seg_22_5_sp4_h_r_7_87262),
    .O(seg_22_7_sp4_v_b_25_83557)
  );
  LocalMux t6474 (
    .I(seg_22_8_sp4_v_b_14_83559),
    .O(seg_22_8_local_g1_6_87542)
  );
  Span4Mux_v3 t6475 (
    .I(seg_22_5_sp4_h_r_9_87264),
    .O(seg_22_8_sp4_v_b_14_83559)
  );
  LocalMux t6476 (
    .I(seg_22_7_sp4_v_b_29_83561),
    .O(seg_22_7_local_g3_5_87434)
  );
  Span4Mux_v2 t6477 (
    .I(seg_22_5_sp4_h_r_11_87256),
    .O(seg_22_7_sp4_v_b_29_83561)
  );
  LocalMux t6478 (
    .I(seg_21_7_sp4_h_r_3_83673),
    .O(seg_21_7_local_g0_3_83577)
  );
  Span4Mux_h4 t6479 (
    .I(seg_25_7_sp4_v_b_10_94851),
    .O(seg_21_7_sp4_h_r_3_83673)
  );
  CascadeMux t648 (
    .I(net_49009),
    .O(net_49009_cascademuxed)
  );
  LocalMux t6480 (
    .I(seg_20_5_sp4_r_v_b_23_79368),
    .O(seg_20_5_local_g3_7_79528)
  );
  Span4Mux_v1 t6481 (
    .I(seg_21_6_sp4_h_r_10_83547),
    .O(seg_20_5_sp4_r_v_b_23_79368)
  );
  Span4Mux_h4 t6482 (
    .I(seg_25_6_sp4_h_r_10_99458),
    .O(seg_21_6_sp4_h_r_10_83547)
  );
  LocalMux t6483 (
    .I(seg_20_5_sp4_v_b_12_76093),
    .O(seg_20_5_local_g0_4_79501)
  );
  Span4Mux_v1 t6484 (
    .I(seg_20_6_sp4_h_r_1_79715),
    .O(seg_20_5_sp4_v_b_12_76093)
  );
  Span4Mux_h4 t6485 (
    .I(seg_24_6_sp4_h_r_1_95107),
    .O(seg_20_6_sp4_h_r_1_79715)
  );
  LocalMux t6486 (
    .I(seg_20_5_sp4_v_b_15_76096),
    .O(seg_20_5_local_g0_7_79504)
  );
  Span4Mux_v1 t6487 (
    .I(seg_20_6_sp4_h_r_2_79718),
    .O(seg_20_5_sp4_v_b_15_76096)
  );
  Span4Mux_h4 t6488 (
    .I(seg_24_6_sp4_h_r_11_95109),
    .O(seg_20_6_sp4_h_r_2_79718)
  );
  LocalMux t6489 (
    .I(seg_23_9_sp4_v_b_21_87520),
    .O(seg_23_9_local_g1_5_91495)
  );
  CascadeMux t649 (
    .I(net_49148),
    .O(net_49148_cascademuxed)
  );
  Span4Mux_v3 t6490 (
    .I(seg_23_6_sp4_h_r_8_91217),
    .O(seg_23_9_sp4_v_b_21_87520)
  );
  LocalMux t6491 (
    .I(seg_22_9_sp4_r_v_b_23_87522),
    .O(seg_22_9_local_g3_7_87682)
  );
  Span4Mux_v3 t6492 (
    .I(seg_23_6_sp4_h_r_10_91209),
    .O(seg_22_9_sp4_r_v_b_23_87522)
  );
  LocalMux t6493 (
    .I(seg_21_9_sp4_r_v_b_12_83680),
    .O(seg_21_9_local_g2_4_83840)
  );
  Span4Mux_v3 t6494 (
    .I(seg_22_6_sp4_h_r_1_87377),
    .O(seg_21_9_sp4_r_v_b_12_83680)
  );
  LocalMux t6495 (
    .I(seg_17_3_sp4_r_v_b_36_68495),
    .O(seg_17_3_local_g2_4_68409)
  );
  Span4Mux_v3 t6496 (
    .I(seg_18_6_sp4_h_r_1_72684),
    .O(seg_17_3_sp4_r_v_b_36_68495)
  );
  Span4Mux_h4 t6497 (
    .I(seg_22_6_sp4_h_r_5_87383),
    .O(seg_18_6_sp4_h_r_1_72684)
  );
  LocalMux t6498 (
    .I(seg_21_4_sp4_h_r_6_83307),
    .O(seg_21_4_local_g1_6_83219)
  );
  Span4Mux_h4 t6499 (
    .I(seg_25_4_sp4_v_t_43_94986),
    .O(seg_21_4_sp4_h_r_6_83307)
  );
  CascadeMux t65 (
    .I(net_11499),
    .O(net_11499_cascademuxed)
  );
  LocalMux t6500 (
    .I(seg_23_5_sp4_v_b_24_87143),
    .O(seg_23_5_local_g3_0_91014)
  );
  Span4Mux_v2 t6501 (
    .I(seg_23_7_sp4_h_r_0_91330),
    .O(seg_23_5_sp4_v_b_24_87143)
  );
  LocalMux t6502 (
    .I(seg_21_5_sp4_r_v_b_24_83312),
    .O(seg_21_5_local_g0_0_83328)
  );
  Span4Mux_v2 t6503 (
    .I(seg_22_7_sp4_h_r_7_87508),
    .O(seg_21_5_sp4_r_v_b_24_83312)
  );
  LocalMux t6504 (
    .I(seg_22_5_sp4_v_b_26_83314),
    .O(seg_22_5_local_g2_2_87177)
  );
  Span4Mux_v2 t6505 (
    .I(seg_22_7_sp4_h_r_9_87510),
    .O(seg_22_5_sp4_v_b_26_83314)
  );
  LocalMux t6506 (
    .I(seg_22_3_sp4_h_r_11_87010),
    .O(seg_22_3_local_g1_3_86924)
  );
  Span4Mux_h0 t6507 (
    .I(seg_22_3_sp4_v_t_46_83321),
    .O(seg_22_3_sp4_h_r_11_87010)
  );
  Span4Mux_v4 t6508 (
    .I(seg_22_7_sp4_h_r_11_87502),
    .O(seg_22_3_sp4_v_t_46_83321)
  );
  LocalMux t6509 (
    .I(seg_20_3_sp4_r_v_b_11_79104),
    .O(seg_20_3_local_g2_3_79270)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t651 (
    .carryinitin(),
    .carryinitout(t650)
  );
  Span4Mux_v1 t6510 (
    .I(seg_21_3_sp4_h_r_6_83184),
    .O(seg_20_3_sp4_r_v_b_11_79104)
  );
  Span4Mux_h4 t6511 (
    .I(seg_25_3_sp4_v_t_37_94841),
    .O(seg_21_3_sp4_h_r_6_83184)
  );
  LocalMux t6512 (
    .I(seg_17_3_sp4_h_r_10_68485),
    .O(seg_17_3_local_g0_2_68391)
  );
  Span4Mux_h4 t6513 (
    .I(seg_21_3_sp4_h_r_2_83180),
    .O(seg_17_3_sp4_h_r_10_68485)
  );
  Span4Mux_h4 t6514 (
    .I(seg_25_3_sp4_v_t_39_94843),
    .O(seg_21_3_sp4_h_r_2_83180)
  );
  LocalMux t6515 (
    .I(seg_15_4_sp4_h_r_30_53292),
    .O(seg_15_4_local_g3_6_60880)
  );
  Span4Mux_h2 t6516 (
    .I(seg_17_4_sp4_h_r_3_68611),
    .O(seg_15_4_sp4_h_r_30_53292)
  );
  Span4Mux_h4 t6517 (
    .I(seg_21_4_sp4_h_r_3_83304),
    .O(seg_17_4_sp4_h_r_3_68611)
  );
  Span4Mux_h4 t6518 (
    .I(seg_25_4_sp4_v_t_44_94987),
    .O(seg_21_4_sp4_h_r_3_83304)
  );
  LocalMux t6519 (
    .I(seg_20_5_sp4_r_v_b_14_79359),
    .O(seg_20_5_local_g2_6_79519)
  );
  CascadeMux t652 (
    .I(net_49271),
    .O(net_49271_cascademuxed)
  );
  Span4Mux_v1 t6520 (
    .I(seg_21_6_sp4_h_r_3_83550),
    .O(seg_20_5_sp4_r_v_b_14_79359)
  );
  Span4Mux_h4 t6521 (
    .I(seg_25_6_sp4_v_t_38_95259),
    .O(seg_21_6_sp4_h_r_3_83550)
  );
  LocalMux t6522 (
    .I(seg_23_5_sp4_v_b_36_87265),
    .O(seg_23_5_local_g3_4_91018)
  );
  Span4Mux_v3 t6523 (
    .I(seg_23_8_sp4_h_r_8_91463),
    .O(seg_23_5_sp4_v_b_36_87265)
  );
  LocalMux t6524 (
    .I(seg_21_3_sp4_r_v_b_12_82936),
    .O(seg_21_3_local_g2_4_83102)
  );
  Span4Mux_v1 t6525 (
    .I(seg_22_4_sp4_v_t_40_83438),
    .O(seg_21_3_sp4_r_v_b_12_82936)
  );
  Span4Mux_v4 t6526 (
    .I(seg_22_8_sp4_h_r_5_87629),
    .O(seg_22_4_sp4_v_t_40_83438)
  );
  LocalMux t6527 (
    .I(seg_22_4_sp4_h_r_0_87130),
    .O(seg_22_4_local_g0_0_87036)
  );
  Span4Mux_h0 t6528 (
    .I(seg_22_4_sp4_v_t_42_83440),
    .O(seg_22_4_sp4_h_r_0_87130)
  );
  Span4Mux_v4 t6529 (
    .I(seg_22_8_sp4_h_r_7_87631),
    .O(seg_22_4_sp4_v_t_42_83440)
  );
  LocalMux t6530 (
    .I(seg_22_3_sp4_v_b_20_82945),
    .O(seg_22_3_local_g0_4_86917)
  );
  Span4Mux_v1 t6531 (
    .I(seg_22_4_sp4_v_t_44_83442),
    .O(seg_22_3_sp4_v_b_20_82945)
  );
  Span4Mux_v4 t6532 (
    .I(seg_22_8_sp4_h_r_9_87633),
    .O(seg_22_4_sp4_v_t_44_83442)
  );
  LocalMux t6533 (
    .I(seg_20_3_sp4_r_v_b_25_79234),
    .O(seg_20_3_local_g1_1_79260)
  );
  Span4Mux_v2 t6534 (
    .I(seg_21_5_sp4_h_r_1_83423),
    .O(seg_20_3_sp4_r_v_b_25_79234)
  );
  Span4Mux_h4 t6535 (
    .I(seg_25_5_sp4_v_t_42_95124),
    .O(seg_21_5_sp4_h_r_1_83423)
  );
  LocalMux t6536 (
    .I(seg_23_5_sp4_h_r_35_83425),
    .O(seg_23_5_local_g2_3_91009)
  );
  Span4Mux_h2 t6537 (
    .I(seg_25_5_sp4_v_t_46_95128),
    .O(seg_23_5_sp4_h_r_35_83425)
  );
  LocalMux t6538 (
    .I(seg_20_5_sp4_r_v_b_22_79367),
    .O(seg_20_5_local_g3_6_79527)
  );
  Span4Mux_v1 t6539 (
    .I(seg_21_6_sp4_h_r_6_83553),
    .O(seg_20_5_sp4_r_v_b_22_79367)
  );
  Span4Mux_h4 t6540 (
    .I(seg_25_6_sp4_v_t_43_95264),
    .O(seg_21_6_sp4_h_r_6_83553)
  );
  LocalMux t6541 (
    .I(seg_20_3_sp4_r_v_b_20_79114),
    .O(seg_20_3_local_g3_4_79279)
  );
  Span4Mux_v1 t6542 (
    .I(seg_21_4_sp4_h_r_4_83305),
    .O(seg_20_3_sp4_r_v_b_20_79114)
  );
  Span4Mux_h4 t6543 (
    .I(seg_25_4_sp4_v_t_41_94984),
    .O(seg_21_4_sp4_h_r_4_83305)
  );
  LocalMux t6544 (
    .I(seg_23_8_sp4_v_b_29_87515),
    .O(seg_23_8_local_g2_5_91380)
  );
  Span4Mux_v2 t6545 (
    .I(seg_23_10_sp4_h_r_0_91699),
    .O(seg_23_8_sp4_v_b_29_87515)
  );
  LocalMux t6546 (
    .I(seg_22_9_sp4_r_v_b_18_87517),
    .O(seg_22_9_local_g3_2_87677)
  );
  Span4Mux_v1 t6547 (
    .I(seg_23_10_sp4_h_r_2_91703),
    .O(seg_22_9_sp4_r_v_b_18_87517)
  );
  LocalMux t6548 (
    .I(seg_22_9_sp4_r_v_b_17_87516),
    .O(seg_22_9_local_g3_1_87676)
  );
  Span4Mux_v1 t6549 (
    .I(seg_23_10_sp4_h_r_4_91705),
    .O(seg_22_9_sp4_r_v_b_17_87516)
  );
  LocalMux t6550 (
    .I(seg_22_8_sp4_r_v_b_27_87513),
    .O(seg_22_8_local_g1_3_87539)
  );
  Span4Mux_v2 t6551 (
    .I(seg_23_10_sp4_h_r_10_91701),
    .O(seg_22_8_sp4_r_v_b_27_87513)
  );
  LocalMux t6552 (
    .I(seg_22_8_sp4_v_b_30_83687),
    .O(seg_22_8_local_g2_6_87550)
  );
  Span4Mux_v2 t6553 (
    .I(seg_22_10_sp4_h_r_1_87869),
    .O(seg_22_8_sp4_v_b_30_83687)
  );
  LocalMux t6554 (
    .I(seg_22_9_sp4_v_b_14_83682),
    .O(seg_22_9_local_g1_6_87665)
  );
  Span4Mux_v1 t6555 (
    .I(seg_22_10_sp4_h_r_3_87873),
    .O(seg_22_9_sp4_v_b_14_83682)
  );
  LocalMux t6556 (
    .I(seg_22_8_sp4_v_b_35_83690),
    .O(seg_22_8_local_g2_3_87547)
  );
  Span4Mux_v2 t6557 (
    .I(seg_22_10_sp4_h_r_11_87871),
    .O(seg_22_8_sp4_v_b_35_83690)
  );
  LocalMux t6558 (
    .I(seg_21_9_sp4_v_b_23_79860),
    .O(seg_21_9_local_g1_7_83835)
  );
  Span4Mux_v1 t6559 (
    .I(seg_21_10_sp4_h_r_5_84044),
    .O(seg_21_9_sp4_v_b_23_79860)
  );
  CascadeMux t656 (
    .I(net_49289),
    .O(net_49289_cascademuxed)
  );
  Span4Mux_h4 t6560 (
    .I(seg_25_10_sp4_v_b_0_95258),
    .O(seg_21_10_sp4_h_r_5_84044)
  );
  LocalMux t6561 (
    .I(seg_21_10_sp4_v_b_15_79975),
    .O(seg_21_10_local_g1_7_83958)
  );
  Span4Mux_v1 t6562 (
    .I(seg_21_11_sp4_h_r_2_84164),
    .O(seg_21_10_sp4_v_b_15_79975)
  );
  Span4Mux_h4 t6563 (
    .I(seg_25_11_sp4_h_r_2_100240),
    .O(seg_21_11_sp4_h_r_2_84164)
  );
  LocalMux t6564 (
    .I(seg_22_9_sp4_v_b_25_83803),
    .O(seg_22_9_local_g2_1_87668)
  );
  Span4Mux_v2 t6565 (
    .I(seg_22_11_sp4_h_r_1_87992),
    .O(seg_22_9_sp4_v_b_25_83803)
  );
  LocalMux t6566 (
    .I(seg_22_4_sp4_v_b_42_83317),
    .O(seg_22_4_local_g2_2_87054)
  );
  Span4Mux_v3 t6567 (
    .I(seg_22_7_sp4_v_t_41_83808),
    .O(seg_22_4_sp4_v_b_42_83317)
  );
  Span4Mux_v4 t6568 (
    .I(seg_22_11_sp4_h_r_11_87994),
    .O(seg_22_7_sp4_v_t_41_83808)
  );
  LocalMux t6569 (
    .I(seg_21_10_sp4_v_b_19_79979),
    .O(seg_21_10_local_g1_3_83954)
  );
  CascadeMux t657 (
    .I(net_49295),
    .O(net_49295_cascademuxed)
  );
  Span4Mux_v3 t6570 (
    .I(seg_21_7_sp4_h_r_0_83668),
    .O(seg_21_10_sp4_v_b_19_79979)
  );
  Span4Mux_h4 t6571 (
    .I(seg_25_7_sp4_v_t_37_95397),
    .O(seg_21_7_sp4_h_r_0_83668)
  );
  LocalMux t6572 (
    .I(seg_20_5_sp4_r_v_b_27_79482),
    .O(seg_20_5_local_g1_3_79508)
  );
  Span4Mux_v2 t6573 (
    .I(seg_21_7_sp4_h_r_10_83670),
    .O(seg_20_5_sp4_r_v_b_27_79482)
  );
  Span4Mux_h4 t6574 (
    .I(seg_25_7_sp4_v_t_47_95407),
    .O(seg_21_7_sp4_h_r_10_83670)
  );
  LocalMux t6575 (
    .I(seg_21_4_sp4_h_r_1_83300),
    .O(seg_21_4_local_g0_1_83206)
  );
  Span4Mux_h4 t6576 (
    .I(seg_25_4_sp4_v_t_36_94979),
    .O(seg_21_4_sp4_h_r_1_83300)
  );
  Span4Mux_v4 t6577 (
    .I(seg_25_8_sp4_v_t_36_95535),
    .O(seg_25_4_sp4_v_t_36_94979)
  );
  LocalMux t6578 (
    .I(seg_18_8_sp4_h_r_21_69108),
    .O(seg_18_8_local_g0_5_72840)
  );
  Span4Mux_h3 t6579 (
    .I(seg_21_8_sp4_h_r_5_83798),
    .O(seg_18_8_sp4_h_r_21_69108)
  );
  CascadeMux t658 (
    .I(net_49400),
    .O(net_49400_cascademuxed)
  );
  Span4Mux_h4 t6580 (
    .I(seg_25_8_sp4_v_t_46_95545),
    .O(seg_21_8_sp4_h_r_5_83798)
  );
  LocalMux t6581 (
    .I(seg_21_4_sp4_v_b_39_79483),
    .O(seg_21_4_local_g3_7_83236)
  );
  Span4Mux_v3 t6582 (
    .I(seg_21_7_sp4_h_r_2_83672),
    .O(seg_21_4_sp4_v_b_39_79483)
  );
  Span4Mux_h4 t6583 (
    .I(seg_25_7_sp4_v_t_45_95405),
    .O(seg_21_7_sp4_h_r_2_83672)
  );
  LocalMux t6584 (
    .I(seg_23_6_sp4_v_b_28_87270),
    .O(seg_23_6_local_g2_4_91133)
  );
  Span4Mux_v2 t6585 (
    .I(seg_23_8_sp4_v_t_41_87762),
    .O(seg_23_6_sp4_v_b_28_87270)
  );
  Span4Mux_v4 t6586 (
    .I(seg_23_12_sp4_h_r_4_91951),
    .O(seg_23_8_sp4_v_t_41_87762)
  );
  LocalMux t6587 (
    .I(seg_21_6_sp4_r_v_b_25_83434),
    .O(seg_21_6_local_g0_1_83452)
  );
  Span4Mux_v2 t6588 (
    .I(seg_22_8_sp4_v_t_40_83930),
    .O(seg_21_6_sp4_r_v_b_25_83434)
  );
  Span4Mux_v4 t6589 (
    .I(seg_22_12_sp4_h_r_5_88121),
    .O(seg_22_8_sp4_v_t_40_83930)
  );
  CascadeMux t659 (
    .I(net_49418),
    .O(net_49418_cascademuxed)
  );
  LocalMux t6590 (
    .I(seg_18_6_sp4_v_b_31_68747),
    .O(seg_18_6_local_g2_7_72612)
  );
  Span4Mux_v2 t6591 (
    .I(seg_18_8_sp4_v_t_46_69243),
    .O(seg_18_6_sp4_v_b_31_68747)
  );
  Span4Mux_v4 t6592 (
    .I(seg_18_12_sp4_h_r_11_73424),
    .O(seg_18_8_sp4_v_t_46_69243)
  );
  Span4Mux_h4 t6593 (
    .I(seg_22_12_sp4_h_r_11_88117),
    .O(seg_18_12_sp4_h_r_11_73424)
  );
  LocalMux t6594 (
    .I(seg_20_5_sp4_r_v_b_41_79608),
    .O(seg_20_5_local_g3_1_79522)
  );
  Span4Mux_v3 t6595 (
    .I(seg_21_8_sp4_h_r_4_83797),
    .O(seg_20_5_sp4_r_v_b_41_79608)
  );
  Span4Mux_h4 t6596 (
    .I(seg_25_8_sp4_v_t_47_95546),
    .O(seg_21_8_sp4_h_r_4_83797)
  );
  LocalMux t6597 (
    .I(seg_17_9_sp4_h_r_1_69222),
    .O(seg_17_9_local_g0_1_69128)
  );
  Span4Mux_h4 t6598 (
    .I(seg_21_9_sp4_h_r_5_83921),
    .O(seg_17_9_sp4_h_r_1_69222)
  );
  Span4Mux_h4 t6599 (
    .I(seg_25_9_sp4_v_t_40_95678),
    .O(seg_21_9_sp4_h_r_5_83921)
  );
  CascadeMux t66 (
    .I(net_11505),
    .O(net_11505_cascademuxed)
  );
  CascadeMux t660 (
    .I(net_49430),
    .O(net_49430_cascademuxed)
  );
  LocalMux t6600 (
    .I(seg_21_5_sp4_v_b_45_79612),
    .O(seg_21_5_local_g3_5_83357)
  );
  Span4Mux_v3 t6601 (
    .I(seg_21_8_sp4_h_r_8_83801),
    .O(seg_21_5_sp4_v_b_45_79612)
  );
  Span4Mux_h4 t6602 (
    .I(seg_25_8_sp4_v_t_39_95538),
    .O(seg_21_8_sp4_h_r_8_83801)
  );
  LocalMux t6603 (
    .I(seg_16_9_sp4_r_v_b_6_65040),
    .O(seg_16_9_local_g1_6_65310)
  );
  Span4Mux_v1 t6604 (
    .I(seg_17_9_sp4_h_r_6_69229),
    .O(seg_16_9_sp4_r_v_b_6_65040)
  );
  Span4Mux_h4 t6605 (
    .I(seg_21_9_sp4_h_r_3_83919),
    .O(seg_17_9_sp4_h_r_6_69229)
  );
  Span4Mux_h4 t6606 (
    .I(seg_25_9_sp4_v_t_44_95682),
    .O(seg_21_9_sp4_h_r_3_83919)
  );
  LocalMux t6607 (
    .I(seg_21_7_sp4_v_b_13_79604),
    .O(seg_21_7_local_g0_5_83579)
  );
  Span4Mux_v1 t6608 (
    .I(seg_21_8_sp4_h_r_0_83791),
    .O(seg_21_7_sp4_v_b_13_79604)
  );
  Span4Mux_h4 t6609 (
    .I(seg_25_8_sp4_v_t_43_95542),
    .O(seg_21_8_sp4_h_r_0_83791)
  );
  CascadeMux t661 (
    .I(net_49517),
    .O(net_49517_cascademuxed)
  );
  LocalMux t6610 (
    .I(seg_23_6_sp4_r_v_b_40_91223),
    .O(seg_23_6_local_g3_0_91137)
  );
  Span4Mux_v3 t6611 (
    .I(seg_24_9_sp4_v_t_44_91719),
    .O(seg_23_6_sp4_r_v_b_40_91223)
  );
  Span4Mux_v4 t6612 (
    .I(seg_24_13_sp4_h_r_9_96090),
    .O(seg_24_9_sp4_v_t_44_91719)
  );
  LocalMux t6613 (
    .I(seg_23_6_sp4_v_b_44_87396),
    .O(seg_23_6_local_g3_4_91141)
  );
  Span4Mux_v3 t6614 (
    .I(seg_23_9_sp4_v_t_43_87887),
    .O(seg_23_6_sp4_v_b_44_87396)
  );
  Span4Mux_v4 t6615 (
    .I(seg_23_13_sp4_h_r_6_92076),
    .O(seg_23_9_sp4_v_t_43_87887)
  );
  LocalMux t6616 (
    .I(seg_22_3_sp4_v_b_35_83075),
    .O(seg_22_3_local_g3_3_86940)
  );
  Span4Mux_v2 t6617 (
    .I(seg_22_5_sp4_v_t_46_83567),
    .O(seg_22_3_sp4_v_b_35_83075)
  );
  Span4Mux_v4 t6618 (
    .I(seg_22_9_sp4_v_t_45_84058),
    .O(seg_22_5_sp4_v_t_46_83567)
  );
  Span4Mux_v4 t6619 (
    .I(seg_22_13_sp4_h_r_3_88242),
    .O(seg_22_9_sp4_v_t_45_84058)
  );
  CascadeMux t662 (
    .I(net_49640),
    .O(net_49640_cascademuxed)
  );
  LocalMux t6620 (
    .I(seg_22_6_sp4_v_b_43_83564),
    .O(seg_22_6_local_g2_3_87301)
  );
  Span4Mux_v3 t6621 (
    .I(seg_22_9_sp4_v_t_47_84060),
    .O(seg_22_6_sp4_v_b_43_83564)
  );
  Span4Mux_v4 t6622 (
    .I(seg_22_13_sp4_h_r_5_88244),
    .O(seg_22_9_sp4_v_t_47_84060)
  );
  LocalMux t6623 (
    .I(seg_22_8_sp4_v_b_15_83560),
    .O(seg_22_8_local_g1_7_87543)
  );
  Span4Mux_v1 t6624 (
    .I(seg_22_9_sp4_v_t_39_84052),
    .O(seg_22_8_sp4_v_b_15_83560)
  );
  Span4Mux_v4 t6625 (
    .I(seg_22_13_sp4_h_r_9_88248),
    .O(seg_22_9_sp4_v_t_39_84052)
  );
  LocalMux t6626 (
    .I(seg_22_5_sp4_h_r_20_83433),
    .O(seg_22_5_local_g0_4_87163)
  );
  Span4Mux_h3 t6627 (
    .I(seg_25_5_sp4_v_t_38_95120),
    .O(seg_22_5_sp4_h_r_20_83433)
  );
  Span4Mux_v4 t6628 (
    .I(seg_25_9_sp4_v_t_37_95675),
    .O(seg_25_5_sp4_v_t_38_95120)
  );
  LocalMux t6629 (
    .I(seg_23_5_sp4_h_r_31_83431),
    .O(seg_23_5_local_g3_7_91021)
  );
  CascadeMux t663 (
    .I(net_49670),
    .O(net_49670_cascademuxed)
  );
  Span4Mux_h2 t6630 (
    .I(seg_25_5_sp4_v_t_36_95118),
    .O(seg_23_5_sp4_h_r_31_83431)
  );
  Span4Mux_v4 t6631 (
    .I(seg_25_9_sp4_v_t_47_95685),
    .O(seg_25_5_sp4_v_t_36_95118)
  );
  LocalMux t6632 (
    .I(seg_21_6_sp4_v_b_36_79726),
    .O(seg_21_6_local_g2_4_83471)
  );
  Span4Mux_v3 t6633 (
    .I(seg_21_9_sp4_h_r_8_83924),
    .O(seg_21_6_sp4_v_b_36_79726)
  );
  Span4Mux_h4 t6634 (
    .I(seg_25_9_sp4_v_t_39_95677),
    .O(seg_21_9_sp4_h_r_8_83924)
  );
  CascadeMux t664 (
    .I(net_49763),
    .O(net_49763_cascademuxed)
  );
  CascadeMux t665 (
    .I(net_49781),
    .O(net_49781_cascademuxed)
  );
  CascadeMux t666 (
    .I(net_49886),
    .O(net_49886_cascademuxed)
  );
  CascadeMux t667 (
    .I(net_49916),
    .O(net_49916_cascademuxed)
  );
  CascadeMux t668 (
    .I(net_50168),
    .O(net_50168_cascademuxed)
  );
  CascadeMux t669 (
    .I(net_50174),
    .O(net_50174_cascademuxed)
  );
  CascadeMux t67 (
    .I(net_11511),
    .O(net_11511_cascademuxed)
  );
  CascadeMux t670 (
    .I(net_50279),
    .O(net_50279_cascademuxed)
  );
  CascadeMux t671 (
    .I(net_50285),
    .O(net_50285_cascademuxed)
  );
  CascadeMux t672 (
    .I(net_50291),
    .O(net_50291_cascademuxed)
  );
  CascadeMux t673 (
    .I(net_50396),
    .O(net_50396_cascademuxed)
  );
  CascadeMux t674 (
    .I(net_50501),
    .O(net_50501_cascademuxed)
  );
  CascadeMux t675 (
    .I(net_50624),
    .O(net_50624_cascademuxed)
  );
  CascadeMux t676 (
    .I(net_50630),
    .O(net_50630_cascademuxed)
  );
  CascadeMux t677 (
    .I(net_50642),
    .O(net_50642_cascademuxed)
  );
  CascadeMux t678 (
    .I(net_50648),
    .O(net_50648_cascademuxed)
  );
  CascadeMux t679 (
    .I(net_50654),
    .O(net_50654_cascademuxed)
  );
  CascadeMux t68 (
    .I(net_11598),
    .O(net_11598_cascademuxed)
  );
  CascadeMux t680 (
    .I(net_50753),
    .O(net_50753_cascademuxed)
  );
  CascadeMux t681 (
    .I(net_50759),
    .O(net_50759_cascademuxed)
  );
  CascadeMux t682 (
    .I(net_50765),
    .O(net_50765_cascademuxed)
  );
  CascadeMux t683 (
    .I(net_50771),
    .O(net_50771_cascademuxed)
  );
  CascadeMux t684 (
    .I(net_50777),
    .O(net_50777_cascademuxed)
  );
  CascadeMux t685 (
    .I(net_50789),
    .O(net_50789_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t687 (
    .carryinitin(),
    .carryinitout(t686)
  );
  CascadeMux t689 (
    .I(net_50870),
    .O(net_50870_cascademuxed)
  );
  CascadeMux t69 (
    .I(net_11616),
    .O(net_11616_cascademuxed)
  );
  CascadeMux t690 (
    .I(net_50876),
    .O(net_50876_cascademuxed)
  );
  CascadeMux t691 (
    .I(net_50882),
    .O(net_50882_cascademuxed)
  );
  CascadeMux t692 (
    .I(net_50888),
    .O(net_50888_cascademuxed)
  );
  CascadeMux t693 (
    .I(net_50894),
    .O(net_50894_cascademuxed)
  );
  CascadeMux t694 (
    .I(net_50900),
    .O(net_50900_cascademuxed)
  );
  CascadeMux t695 (
    .I(net_50906),
    .O(net_50906_cascademuxed)
  );
  CascadeMux t696 (
    .I(net_50912),
    .O(net_50912_cascademuxed)
  );
  CascadeMux t697 (
    .I(net_50993),
    .O(net_50993_cascademuxed)
  );
  CascadeMux t698 (
    .I(net_50999),
    .O(net_50999_cascademuxed)
  );
  CascadeMux t699 (
    .I(net_51011),
    .O(net_51011_cascademuxed)
  );
  CascadeMux t7 (
    .I(net_6937),
    .O(net_6937_cascademuxed)
  );
  CascadeMux t70 (
    .I(net_11622),
    .O(net_11622_cascademuxed)
  );
  CascadeMux t700 (
    .I(net_51035),
    .O(net_51035_cascademuxed)
  );
  CascadeMux t701 (
    .I(net_52846),
    .O(net_52846_cascademuxed)
  );
  CascadeMux t702 (
    .I(net_52852),
    .O(net_52852_cascademuxed)
  );
  CascadeMux t703 (
    .I(net_52985),
    .O(net_52985_cascademuxed)
  );
  CascadeMux t704 (
    .I(net_53126),
    .O(net_53126_cascademuxed)
  );
  CascadeMux t705 (
    .I(net_53132),
    .O(net_53132_cascademuxed)
  );
  CascadeMux t706 (
    .I(net_53138),
    .O(net_53138_cascademuxed)
  );
  CascadeMux t707 (
    .I(net_53144),
    .O(net_53144_cascademuxed)
  );
  CascadeMux t708 (
    .I(net_53231),
    .O(net_53231_cascademuxed)
  );
  CascadeMux t709 (
    .I(net_53261),
    .O(net_53261_cascademuxed)
  );
  CascadeMux t71 (
    .I(net_11628),
    .O(net_11628_cascademuxed)
  );
  CascadeMux t710 (
    .I(net_53354),
    .O(net_53354_cascademuxed)
  );
  CascadeMux t711 (
    .I(net_53384),
    .O(net_53384_cascademuxed)
  );
  CascadeMux t712 (
    .I(net_53495),
    .O(net_53495_cascademuxed)
  );
  CascadeMux t713 (
    .I(net_53600),
    .O(net_53600_cascademuxed)
  );
  CascadeMux t714 (
    .I(net_53606),
    .O(net_53606_cascademuxed)
  );
  CascadeMux t715 (
    .I(net_53624),
    .O(net_53624_cascademuxed)
  );
  CascadeMux t716 (
    .I(net_53630),
    .O(net_53630_cascademuxed)
  );
  CascadeMux t717 (
    .I(net_53636),
    .O(net_53636_cascademuxed)
  );
  CascadeMux t718 (
    .I(net_53717),
    .O(net_53717_cascademuxed)
  );
  CascadeMux t719 (
    .I(net_53723),
    .O(net_53723_cascademuxed)
  );
  CascadeMux t72 (
    .I(net_11634),
    .O(net_11634_cascademuxed)
  );
  CascadeMux t720 (
    .I(net_53729),
    .O(net_53729_cascademuxed)
  );
  CascadeMux t721 (
    .I(net_53741),
    .O(net_53741_cascademuxed)
  );
  CascadeMux t722 (
    .I(net_53747),
    .O(net_53747_cascademuxed)
  );
  CascadeMux t723 (
    .I(net_53753),
    .O(net_53753_cascademuxed)
  );
  CascadeMux t724 (
    .I(net_53852),
    .O(net_53852_cascademuxed)
  );
  CascadeMux t725 (
    .I(net_53963),
    .O(net_53963_cascademuxed)
  );
  CascadeMux t726 (
    .I(net_53969),
    .O(net_53969_cascademuxed)
  );
  CascadeMux t727 (
    .I(net_53987),
    .O(net_53987_cascademuxed)
  );
  CascadeMux t728 (
    .I(net_54110),
    .O(net_54110_cascademuxed)
  );
  CascadeMux t729 (
    .I(net_54116),
    .O(net_54116_cascademuxed)
  );
  CascadeMux t73 (
    .I(net_11715),
    .O(net_11715_cascademuxed)
  );
  CascadeMux t730 (
    .I(net_54122),
    .O(net_54122_cascademuxed)
  );
  CascadeMux t731 (
    .I(net_54245),
    .O(net_54245_cascademuxed)
  );
  CascadeMux t732 (
    .I(net_54251),
    .O(net_54251_cascademuxed)
  );
  CascadeMux t733 (
    .I(net_54338),
    .O(net_54338_cascademuxed)
  );
  CascadeMux t734 (
    .I(net_54356),
    .O(net_54356_cascademuxed)
  );
  CascadeMux t735 (
    .I(net_54368),
    .O(net_54368_cascademuxed)
  );
  CascadeMux t736 (
    .I(net_54374),
    .O(net_54374_cascademuxed)
  );
  CascadeMux t737 (
    .I(net_54461),
    .O(net_54461_cascademuxed)
  );
  CascadeMux t738 (
    .I(net_54491),
    .O(net_54491_cascademuxed)
  );
  CascadeMux t739 (
    .I(net_54497),
    .O(net_54497_cascademuxed)
  );
  CascadeMux t74 (
    .I(net_11733),
    .O(net_11733_cascademuxed)
  );
  CascadeMux t740 (
    .I(net_54578),
    .O(net_54578_cascademuxed)
  );
  CascadeMux t741 (
    .I(net_54584),
    .O(net_54584_cascademuxed)
  );
  CascadeMux t742 (
    .I(net_54590),
    .O(net_54590_cascademuxed)
  );
  CascadeMux t743 (
    .I(net_54620),
    .O(net_54620_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t745 (
    .carryinitin(),
    .carryinitout(t744)
  );
  CascadeMux t747 (
    .I(net_54707),
    .O(net_54707_cascademuxed)
  );
  CascadeMux t748 (
    .I(net_54719),
    .O(net_54719_cascademuxed)
  );
  CascadeMux t749 (
    .I(net_54725),
    .O(net_54725_cascademuxed)
  );
  CascadeMux t75 (
    .I(net_11739),
    .O(net_11739_cascademuxed)
  );
  CascadeMux t750 (
    .I(net_54731),
    .O(net_54731_cascademuxed)
  );
  CascadeMux t751 (
    .I(net_54737),
    .O(net_54737_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t752 (
    .carryinitin(net_58570),
    .carryinitout(net_58614)
  );
  CascadeMux t753 (
    .I(net_54842),
    .O(net_54842_cascademuxed)
  );
  CascadeMux t754 (
    .I(net_54854),
    .O(net_54854_cascademuxed)
  );
  CascadeMux t755 (
    .I(net_54947),
    .O(net_54947_cascademuxed)
  );
  CascadeMux t756 (
    .I(net_54953),
    .O(net_54953_cascademuxed)
  );
  CascadeMux t757 (
    .I(net_54959),
    .O(net_54959_cascademuxed)
  );
  CascadeMux t758 (
    .I(net_54965),
    .O(net_54965_cascademuxed)
  );
  CascadeMux t759 (
    .I(net_54977),
    .O(net_54977_cascademuxed)
  );
  CascadeMux t76 (
    .I(net_11745),
    .O(net_11745_cascademuxed)
  );
  CascadeMux t760 (
    .I(net_54983),
    .O(net_54983_cascademuxed)
  );
  CascadeMux t761 (
    .I(net_54989),
    .O(net_54989_cascademuxed)
  );
  CascadeMux t762 (
    .I(net_55112),
    .O(net_55112_cascademuxed)
  );
  CascadeMux t763 (
    .I(net_56682),
    .O(net_56682_cascademuxed)
  );
  CascadeMux t764 (
    .I(net_56809),
    .O(net_56809_cascademuxed)
  );
  CascadeMux t765 (
    .I(net_56827),
    .O(net_56827_cascademuxed)
  );
  CascadeMux t766 (
    .I(net_56845),
    .O(net_56845_cascademuxed)
  );
  CascadeMux t767 (
    .I(net_57055),
    .O(net_57055_cascademuxed)
  );
  CascadeMux t768 (
    .I(net_57067),
    .O(net_57067_cascademuxed)
  );
  CascadeMux t769 (
    .I(net_57079),
    .O(net_57079_cascademuxed)
  );
  CascadeMux t77 (
    .I(net_11751),
    .O(net_11751_cascademuxed)
  );
  CascadeMux t770 (
    .I(net_57178),
    .O(net_57178_cascademuxed)
  );
  CascadeMux t771 (
    .I(net_57202),
    .O(net_57202_cascademuxed)
  );
  CascadeMux t772 (
    .I(net_57208),
    .O(net_57208_cascademuxed)
  );
  CascadeMux t773 (
    .I(net_57214),
    .O(net_57214_cascademuxed)
  );
  CascadeMux t774 (
    .I(net_57307),
    .O(net_57307_cascademuxed)
  );
  CascadeMux t775 (
    .I(net_57319),
    .O(net_57319_cascademuxed)
  );
  CascadeMux t776 (
    .I(net_57325),
    .O(net_57325_cascademuxed)
  );
  CascadeMux t777 (
    .I(net_57337),
    .O(net_57337_cascademuxed)
  );
  CascadeMux t778 (
    .I(net_57343),
    .O(net_57343_cascademuxed)
  );
  CascadeMux t779 (
    .I(net_57460),
    .O(net_57460_cascademuxed)
  );
  CascadeMux t78 (
    .I(net_11838),
    .O(net_11838_cascademuxed)
  );
  CascadeMux t780 (
    .I(net_57547),
    .O(net_57547_cascademuxed)
  );
  CascadeMux t781 (
    .I(net_57559),
    .O(net_57559_cascademuxed)
  );
  CascadeMux t782 (
    .I(net_57583),
    .O(net_57583_cascademuxed)
  );
  CascadeMux t783 (
    .I(net_57706),
    .O(net_57706_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t785 (
    .carryinitin(),
    .carryinitout(t784)
  );
  CascadeMux t787 (
    .I(net_57799),
    .O(net_57799_cascademuxed)
  );
  CascadeMux t788 (
    .I(net_57817),
    .O(net_57817_cascademuxed)
  );
  CascadeMux t789 (
    .I(net_57835),
    .O(net_57835_cascademuxed)
  );
  CascadeMux t79 (
    .I(net_11850),
    .O(net_11850_cascademuxed)
  );
  CascadeMux t790 (
    .I(net_57934),
    .O(net_57934_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t792 (
    .carryinitin(),
    .carryinitout(t791)
  );
  CascadeMux t793 (
    .I(net_58174),
    .O(net_58174_cascademuxed)
  );
  CascadeMux t794 (
    .I(net_58180),
    .O(net_58180_cascademuxed)
  );
  CascadeMux t795 (
    .I(net_58186),
    .O(net_58186_cascademuxed)
  );
  CascadeMux t796 (
    .I(net_58198),
    .O(net_58198_cascademuxed)
  );
  CascadeMux t797 (
    .I(net_58204),
    .O(net_58204_cascademuxed)
  );
  CascadeMux t798 (
    .I(net_58285),
    .O(net_58285_cascademuxed)
  );
  CascadeMux t799 (
    .I(net_58321),
    .O(net_58321_cascademuxed)
  );
  CascadeMux t8 (
    .I(net_6943),
    .O(net_6943_cascademuxed)
  );
  CascadeMux t80 (
    .I(net_11862),
    .O(net_11862_cascademuxed)
  );
  CascadeMux t800 (
    .I(net_58327),
    .O(net_58327_cascademuxed)
  );
  CascadeMux t801 (
    .I(net_58444),
    .O(net_58444_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t803 (
    .carryinitin(),
    .carryinitout(t802)
  );
  CascadeMux t805 (
    .I(net_58531),
    .O(net_58531_cascademuxed)
  );
  CascadeMux t806 (
    .I(net_58537),
    .O(net_58537_cascademuxed)
  );
  CascadeMux t807 (
    .I(net_58543),
    .O(net_58543_cascademuxed)
  );
  CascadeMux t808 (
    .I(net_58549),
    .O(net_58549_cascademuxed)
  );
  CascadeMux t809 (
    .I(net_58555),
    .O(net_58555_cascademuxed)
  );
  CascadeMux t81 (
    .I(net_11967),
    .O(net_11967_cascademuxed)
  );
  CascadeMux t810 (
    .I(net_58561),
    .O(net_58561_cascademuxed)
  );
  CascadeMux t811 (
    .I(net_58567),
    .O(net_58567_cascademuxed)
  );
  CascadeMux t812 (
    .I(net_58573),
    .O(net_58573_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t813 (
    .carryinitin(net_62400),
    .carryinitout(net_62444)
  );
  CascadeMux t814 (
    .I(net_58654),
    .O(net_58654_cascademuxed)
  );
  CascadeMux t815 (
    .I(net_58672),
    .O(net_58672_cascademuxed)
  );
  CascadeMux t816 (
    .I(net_58690),
    .O(net_58690_cascademuxed)
  );
  CascadeMux t817 (
    .I(net_58777),
    .O(net_58777_cascademuxed)
  );
  CascadeMux t818 (
    .I(net_58783),
    .O(net_58783_cascademuxed)
  );
  CascadeMux t819 (
    .I(net_58789),
    .O(net_58789_cascademuxed)
  );
  CascadeMux t82 (
    .I(net_11973),
    .O(net_11973_cascademuxed)
  );
  CascadeMux t820 (
    .I(net_58795),
    .O(net_58795_cascademuxed)
  );
  CascadeMux t821 (
    .I(net_58807),
    .O(net_58807_cascademuxed)
  );
  CascadeMux t822 (
    .I(net_58813),
    .O(net_58813_cascademuxed)
  );
  CascadeMux t823 (
    .I(net_58819),
    .O(net_58819_cascademuxed)
  );
  CascadeMux t824 (
    .I(net_58918),
    .O(net_58918_cascademuxed)
  );
  CascadeMux t825 (
    .I(net_60774),
    .O(net_60774_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t827 (
    .carryinitin(),
    .carryinitout(t826)
  );
  CascadeMux t828 (
    .I(net_60909),
    .O(net_60909_cascademuxed)
  );
  CascadeMux t829 (
    .I(net_60915),
    .O(net_60915_cascademuxed)
  );
  CascadeMux t83 (
    .I(net_11979),
    .O(net_11979_cascademuxed)
  );
  CascadeMux t830 (
    .I(net_60921),
    .O(net_60921_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t831 (
    .carryinitin(net_64755),
    .carryinitout(net_64799)
  );
  CascadeMux t832 (
    .I(net_61020),
    .O(net_61020_cascademuxed)
  );
  CascadeMux t833 (
    .I(net_61032),
    .O(net_61032_cascademuxed)
  );
  CascadeMux t834 (
    .I(net_61044),
    .O(net_61044_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t836 (
    .carryinitin(),
    .carryinitout(t835)
  );
  CascadeMux t837 (
    .I(net_61131),
    .O(net_61131_cascademuxed)
  );
  CascadeMux t838 (
    .I(net_61137),
    .O(net_61137_cascademuxed)
  );
  CascadeMux t839 (
    .I(net_61149),
    .O(net_61149_cascademuxed)
  );
  CascadeMux t84 (
    .I(net_11991),
    .O(net_11991_cascademuxed)
  );
  CascadeMux t840 (
    .I(net_61155),
    .O(net_61155_cascademuxed)
  );
  CascadeMux t841 (
    .I(net_61161),
    .O(net_61161_cascademuxed)
  );
  CascadeMux t842 (
    .I(net_61167),
    .O(net_61167_cascademuxed)
  );
  CascadeMux t843 (
    .I(net_61173),
    .O(net_61173_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t844 (
    .carryinitin(net_65001),
    .carryinitout(net_65045)
  );
  CascadeMux t845 (
    .I(net_61266),
    .O(net_61266_cascademuxed)
  );
  CascadeMux t846 (
    .I(net_61272),
    .O(net_61272_cascademuxed)
  );
  CascadeMux t847 (
    .I(net_61290),
    .O(net_61290_cascademuxed)
  );
  CascadeMux t848 (
    .I(net_61395),
    .O(net_61395_cascademuxed)
  );
  CascadeMux t849 (
    .I(net_61506),
    .O(net_61506_cascademuxed)
  );
  CascadeMux t850 (
    .I(net_61524),
    .O(net_61524_cascademuxed)
  );
  CascadeMux t851 (
    .I(net_61536),
    .O(net_61536_cascademuxed)
  );
  CascadeMux t852 (
    .I(net_61641),
    .O(net_61641_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t854 (
    .carryinitin(),
    .carryinitout(t853)
  );
  CascadeMux t855 (
    .I(net_61746),
    .O(net_61746_cascademuxed)
  );
  CascadeMux t856 (
    .I(net_61752),
    .O(net_61752_cascademuxed)
  );
  CascadeMux t857 (
    .I(net_61776),
    .O(net_61776_cascademuxed)
  );
  CascadeMux t858 (
    .I(net_61788),
    .O(net_61788_cascademuxed)
  );
  CascadeMux t859 (
    .I(net_61869),
    .O(net_61869_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t86 (
    .carryinitin(),
    .carryinitout(t85)
  );
  CascadeMux t860 (
    .I(net_61887),
    .O(net_61887_cascademuxed)
  );
  CascadeMux t861 (
    .I(net_61899),
    .O(net_61899_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t863 (
    .carryinitin(),
    .carryinitout(t862)
  );
  CascadeMux t864 (
    .I(net_61992),
    .O(net_61992_cascademuxed)
  );
  CascadeMux t865 (
    .I(net_62004),
    .O(net_62004_cascademuxed)
  );
  CascadeMux t866 (
    .I(net_62010),
    .O(net_62010_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t868 (
    .carryinitin(),
    .carryinitout(t867)
  );
  CascadeMux t869 (
    .I(net_62115),
    .O(net_62115_cascademuxed)
  );
  CascadeMux t87 (
    .I(net_12090),
    .O(net_12090_cascademuxed)
  );
  CascadeMux t870 (
    .I(net_62121),
    .O(net_62121_cascademuxed)
  );
  CascadeMux t871 (
    .I(net_62127),
    .O(net_62127_cascademuxed)
  );
  CascadeMux t872 (
    .I(net_62133),
    .O(net_62133_cascademuxed)
  );
  CascadeMux t873 (
    .I(net_62145),
    .O(net_62145_cascademuxed)
  );
  CascadeMux t874 (
    .I(net_62250),
    .O(net_62250_cascademuxed)
  );
  CascadeMux t875 (
    .I(net_62256),
    .O(net_62256_cascademuxed)
  );
  CascadeMux t876 (
    .I(net_62280),
    .O(net_62280_cascademuxed)
  );
  CascadeMux t877 (
    .I(net_62361),
    .O(net_62361_cascademuxed)
  );
  CascadeMux t878 (
    .I(net_62367),
    .O(net_62367_cascademuxed)
  );
  CascadeMux t879 (
    .I(net_62373),
    .O(net_62373_cascademuxed)
  );
  CascadeMux t88 (
    .I(net_12120),
    .O(net_12120_cascademuxed)
  );
  CascadeMux t880 (
    .I(net_62379),
    .O(net_62379_cascademuxed)
  );
  CascadeMux t881 (
    .I(net_62385),
    .O(net_62385_cascademuxed)
  );
  CascadeMux t882 (
    .I(net_62391),
    .O(net_62391_cascademuxed)
  );
  CascadeMux t883 (
    .I(net_62397),
    .O(net_62397_cascademuxed)
  );
  CascadeMux t884 (
    .I(net_62403),
    .O(net_62403_cascademuxed)
  );
  CascadeMux t885 (
    .I(net_62484),
    .O(net_62484_cascademuxed)
  );
  CascadeMux t886 (
    .I(net_62496),
    .O(net_62496_cascademuxed)
  );
  CascadeMux t887 (
    .I(net_62631),
    .O(net_62631_cascademuxed)
  );
  CascadeMux t888 (
    .I(net_64488),
    .O(net_64488_cascademuxed)
  );
  CascadeMux t889 (
    .I(net_64605),
    .O(net_64605_cascademuxed)
  );
  CascadeMux t89 (
    .I(net_12207),
    .O(net_12207_cascademuxed)
  );
  CascadeMux t890 (
    .I(net_64716),
    .O(net_64716_cascademuxed)
  );
  CascadeMux t891 (
    .I(net_64722),
    .O(net_64722_cascademuxed)
  );
  CascadeMux t892 (
    .I(net_64728),
    .O(net_64728_cascademuxed)
  );
  CascadeMux t893 (
    .I(net_64734),
    .O(net_64734_cascademuxed)
  );
  CascadeMux t894 (
    .I(net_64740),
    .O(net_64740_cascademuxed)
  );
  CascadeMux t895 (
    .I(net_64746),
    .O(net_64746_cascademuxed)
  );
  CascadeMux t896 (
    .I(net_64752),
    .O(net_64752_cascademuxed)
  );
  CascadeMux t897 (
    .I(net_64758),
    .O(net_64758_cascademuxed)
  );
  CascadeMux t898 (
    .I(net_64839),
    .O(net_64839_cascademuxed)
  );
  CascadeMux t899 (
    .I(net_64845),
    .O(net_64845_cascademuxed)
  );
  CascadeMux t9 (
    .I(net_6949),
    .O(net_6949_cascademuxed)
  );
  CascadeMux t90 (
    .I(net_12213),
    .O(net_12213_cascademuxed)
  );
  CascadeMux t900 (
    .I(net_64851),
    .O(net_64851_cascademuxed)
  );
  CascadeMux t901 (
    .I(net_64881),
    .O(net_64881_cascademuxed)
  );
  CascadeMux t902 (
    .I(net_64962),
    .O(net_64962_cascademuxed)
  );
  CascadeMux t903 (
    .I(net_64968),
    .O(net_64968_cascademuxed)
  );
  CascadeMux t904 (
    .I(net_64974),
    .O(net_64974_cascademuxed)
  );
  CascadeMux t905 (
    .I(net_64986),
    .O(net_64986_cascademuxed)
  );
  CascadeMux t906 (
    .I(net_64998),
    .O(net_64998_cascademuxed)
  );
  CascadeMux t907 (
    .I(net_65004),
    .O(net_65004_cascademuxed)
  );
  CascadeMux t908 (
    .I(net_65085),
    .O(net_65085_cascademuxed)
  );
  CascadeMux t909 (
    .I(net_65103),
    .O(net_65103_cascademuxed)
  );
  CascadeMux t91 (
    .I(net_12225),
    .O(net_12225_cascademuxed)
  );
  CascadeMux t910 (
    .I(net_65121),
    .O(net_65121_cascademuxed)
  );
  CascadeMux t911 (
    .I(net_65214),
    .O(net_65214_cascademuxed)
  );
  CascadeMux t912 (
    .I(net_65232),
    .O(net_65232_cascademuxed)
  );
  CascadeMux t913 (
    .I(net_65337),
    .O(net_65337_cascademuxed)
  );
  CascadeMux t914 (
    .I(net_65454),
    .O(net_65454_cascademuxed)
  );
  CascadeMux t915 (
    .I(net_65472),
    .O(net_65472_cascademuxed)
  );
  CascadeMux t916 (
    .I(net_65478),
    .O(net_65478_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t918 (
    .carryinitin(),
    .carryinitout(t917)
  );
  CascadeMux t919 (
    .I(net_65577),
    .O(net_65577_cascademuxed)
  );
  CascadeMux t92 (
    .I(net_12231),
    .O(net_12231_cascademuxed)
  );
  CascadeMux t920 (
    .I(net_65583),
    .O(net_65583_cascademuxed)
  );
  CascadeMux t921 (
    .I(net_65589),
    .O(net_65589_cascademuxed)
  );
  CascadeMux t922 (
    .I(net_65595),
    .O(net_65595_cascademuxed)
  );
  CascadeMux t923 (
    .I(net_65601),
    .O(net_65601_cascademuxed)
  );
  CascadeMux t924 (
    .I(net_65613),
    .O(net_65613_cascademuxed)
  );
  CascadeMux t925 (
    .I(net_65712),
    .O(net_65712_cascademuxed)
  );
  CascadeMux t926 (
    .I(net_65718),
    .O(net_65718_cascademuxed)
  );
  CascadeMux t927 (
    .I(net_65736),
    .O(net_65736_cascademuxed)
  );
  CascadeMux t928 (
    .I(net_65742),
    .O(net_65742_cascademuxed)
  );
  CascadeMux t93 (
    .I(net_12249),
    .O(net_12249_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t930 (
    .carryinitin(),
    .carryinitout(t929)
  );
  CascadeMux t931 (
    .I(net_65823),
    .O(net_65823_cascademuxed)
  );
  CascadeMux t932 (
    .I(net_65829),
    .O(net_65829_cascademuxed)
  );
  CascadeMux t933 (
    .I(net_65835),
    .O(net_65835_cascademuxed)
  );
  CascadeMux t934 (
    .I(net_65841),
    .O(net_65841_cascademuxed)
  );
  CascadeMux t935 (
    .I(net_65847),
    .O(net_65847_cascademuxed)
  );
  CascadeMux t936 (
    .I(net_65853),
    .O(net_65853_cascademuxed)
  );
  CascadeMux t937 (
    .I(net_65946),
    .O(net_65946_cascademuxed)
  );
  CascadeMux t938 (
    .I(net_65952),
    .O(net_65952_cascademuxed)
  );
  CascadeMux t939 (
    .I(net_65958),
    .O(net_65958_cascademuxed)
  );
  CascadeMux t940 (
    .I(net_65964),
    .O(net_65964_cascademuxed)
  );
  CascadeMux t941 (
    .I(net_65970),
    .O(net_65970_cascademuxed)
  );
  CascadeMux t942 (
    .I(net_65976),
    .O(net_65976_cascademuxed)
  );
  CascadeMux t943 (
    .I(net_65982),
    .O(net_65982_cascademuxed)
  );
  CascadeMux t944 (
    .I(net_65988),
    .O(net_65988_cascademuxed)
  );
  CascadeMux t945 (
    .I(net_66069),
    .O(net_66069_cascademuxed)
  );
  CascadeMux t946 (
    .I(net_66075),
    .O(net_66075_cascademuxed)
  );
  CascadeMux t947 (
    .I(net_66105),
    .O(net_66105_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t949 (
    .carryinitin(),
    .carryinitout(t948)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t95 (
    .carryinitin(),
    .carryinitout(t94)
  );
  CascadeMux t950 (
    .I(net_66192),
    .O(net_66192_cascademuxed)
  );
  CascadeMux t951 (
    .I(net_66198),
    .O(net_66198_cascademuxed)
  );
  CascadeMux t952 (
    .I(net_66204),
    .O(net_66204_cascademuxed)
  );
  CascadeMux t953 (
    .I(net_66210),
    .O(net_66210_cascademuxed)
  );
  CascadeMux t954 (
    .I(net_66216),
    .O(net_66216_cascademuxed)
  );
  CascadeMux t955 (
    .I(net_66228),
    .O(net_66228_cascademuxed)
  );
  CascadeMux t956 (
    .I(net_66234),
    .O(net_66234_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t958 (
    .carryinitin(net_70062),
    .carryinitout(net_70106)
  );
  CascadeMux t959 (
    .I(net_66315),
    .O(net_66315_cascademuxed)
  );
  CascadeMux t96 (
    .I(net_12477),
    .O(net_12477_cascademuxed)
  );
  CascadeMux t960 (
    .I(net_66321),
    .O(net_66321_cascademuxed)
  );
  CascadeMux t961 (
    .I(net_66327),
    .O(net_66327_cascademuxed)
  );
  CascadeMux t962 (
    .I(net_66345),
    .O(net_66345_cascademuxed)
  );
  CascadeMux t963 (
    .I(net_66357),
    .O(net_66357_cascademuxed)
  );
  CascadeMux t964 (
    .I(net_66438),
    .O(net_66438_cascademuxed)
  );
  CascadeMux t965 (
    .I(net_68424),
    .O(net_68424_cascademuxed)
  );
  CascadeMux t966 (
    .I(net_68430),
    .O(net_68430_cascademuxed)
  );
  CascadeMux t967 (
    .I(net_68436),
    .O(net_68436_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t969 (
    .carryinitin(),
    .carryinitout(t968)
  );
  CascadeMux t97 (
    .I(net_12483),
    .O(net_12483_cascademuxed)
  );
  CascadeMux t970 (
    .I(net_68553),
    .O(net_68553_cascademuxed)
  );
  CascadeMux t971 (
    .I(net_68583),
    .O(net_68583_cascademuxed)
  );
  CascadeMux t972 (
    .I(net_68589),
    .O(net_68589_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t973 (
    .carryinitin(net_72417),
    .carryinitout(net_72461)
  );
  CascadeMux t974 (
    .I(net_68670),
    .O(net_68670_cascademuxed)
  );
  CascadeMux t975 (
    .I(net_68682),
    .O(net_68682_cascademuxed)
  );
  CascadeMux t976 (
    .I(net_68706),
    .O(net_68706_cascademuxed)
  );
  CascadeMux t977 (
    .I(net_68712),
    .O(net_68712_cascademuxed)
  );
  CascadeMux t978 (
    .I(net_68805),
    .O(net_68805_cascademuxed)
  );
  CascadeMux t979 (
    .I(net_68835),
    .O(net_68835_cascademuxed)
  );
  CascadeMux t98 (
    .I(net_12576),
    .O(net_12576_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t981 (
    .carryinitin(),
    .carryinitout(t980)
  );
  CascadeMux t982 (
    .I(net_68958),
    .O(net_68958_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t983 (
    .carryinitin(net_72786),
    .carryinitout(net_72830)
  );
  CascadeMux t984 (
    .I(net_69045),
    .O(net_69045_cascademuxed)
  );
  CascadeMux t985 (
    .I(net_69051),
    .O(net_69051_cascademuxed)
  );
  CascadeMux t986 (
    .I(net_69075),
    .O(net_69075_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t988 (
    .carryinitin(),
    .carryinitout(t987)
  );
  CascadeMux t989 (
    .I(net_69303),
    .O(net_69303_cascademuxed)
  );
  CascadeMux t99 (
    .I(net_12582),
    .O(net_12582_cascademuxed)
  );
  CascadeMux t990 (
    .I(net_69408),
    .O(net_69408_cascademuxed)
  );
  CascadeMux t991 (
    .I(net_69414),
    .O(net_69414_cascademuxed)
  );
  CascadeMux t992 (
    .I(net_69420),
    .O(net_69420_cascademuxed)
  );
  CascadeMux t993 (
    .I(net_69426),
    .O(net_69426_cascademuxed)
  );
  CascadeMux t994 (
    .I(net_69438),
    .O(net_69438_cascademuxed)
  );
  CascadeMux t995 (
    .I(net_69549),
    .O(net_69549_cascademuxed)
  );
  CascadeMux t996 (
    .I(net_69555),
    .O(net_69555_cascademuxed)
  );
  CascadeMux t997 (
    .I(net_69654),
    .O(net_69654_cascademuxed)
  );
  CascadeMux t998 (
    .I(net_69660),
    .O(net_69660_cascademuxed)
  );
  CascadeMux t999 (
    .I(net_69666),
    .O(net_69666_cascademuxed)
  );
endmodule
