//==============================================================================
// DFT Twiddle Factors ROM
//
// 16-bit twiddle factor formula for N-point window DFT:
//   w_i = int(exp(2 * pi * j * i / N) * (2^15)),
// where
//  i = 0 ... N
//
// However, for enveloppe extraction we need only 3 points: w_1, w_2, w_3.
//
//==============================================================================

module dft_twiddle_rom
#(
    parameter ADDR_W = 2,   // Memory depth
    parameter DATA_W = 16  // Data width
)(
    // System
    input wire               clk,       // System clock
    input wire               rst,       // System reset
    // Read interface
    output wire [DATA_W-1:0] rdata_re, // Read data real part
    output wire [DATA_W-1:0] rdata_im, // Read data imaginary part
    input  wire [ADDR_W-1:0] raddr,    // Read address
    input  wire              rd        // Read enable
);

`ifdef YOSYS
  `define IP_LEGACY
`elsif __ICARUS__
  `define IP_LEGACY
`endif

`ifdef IP_LEGACY
 SB_RAM40_4K #(
    .INIT_0(256'h000000000000000000000000000000000000000000000000000030fc5a827642),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),

    .INIT_FILE("../../rtl/mem_files/dft_twiddle_re_16.mem"),
    .READ_MODE(2'h0),
    .WRITE_MODE(2'h0)
) mem_re (
    .MASK(16'h0000),
    .RADDR({{11-ADDR_W{1'b0}}, raddr}),
    .RCLK(clk),
    .RCLKE(1'h1),
    .RDATA(rdata_re),
    .RE(1'h1),
    .WADDR(11'h000),
    .WCLK(clk),
    .WCLKE(1'h1),
    .WDATA(16'h0000),
    .WE(1'h0)
);

SB_RAM40_4K #(
    .INIT_0(256'h000000000000000000000000000000000000000000000000000076425a8230fc),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),

    .INIT_FILE("../../rtl/mem_files/dft_twiddle_im_16.mem"),
    .READ_MODE(2'h0),
    .WRITE_MODE(2'h0)
) mem_im (
    .MASK(16'h0000),
    .RADDR({{11-ADDR_W{1'b0}}, raddr}),
    .RCLK(clk),
    .RCLKE(1'h1),
    .RDATA(rdata_im),
    .RE(1'h1),
    .WADDR(11'h000),
    .WCLK(clk),
    .WCLKE(1'h1),
    .WDATA(16'h0000),
    .WE(1'h0)
);

`else

PDP4K #(
    .INITVAL_0("0x000000000000000000000000000000000000000000000000000030fc5a827642"),
    .INITVAL_1("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_2("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_3("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_4("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_5("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_6("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_7("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_8("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_9("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_A("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_B("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_C("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_D("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_E("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_F("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .DATA_WIDTH_W("16"),
    .DATA_WIDTH_R("16")
) mem_re (
    .DI     (16'h0000),
    .ADW    (11'h000),
    .ADR    ({{11-ADDR_W{1'b0}}, raddr}),
    .CKW    (clk),
    .CKR    (clk),
    .CEW    (1'h1),
    .CER    (1'h1),
    .RE     (1'h1),
    .WE     (1'h0),
    .MASK_N (16'h0000),
    .DO     (rdata_re)
);

PDP4K #(
    .INITVAL_0("0x000000000000000000000000000000000000000000000000000076425a8230fc"),
    .INITVAL_1("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_2("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_3("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_4("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_5("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_6("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_7("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_8("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_9("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_A("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_B("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_C("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_D("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_E("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .INITVAL_F("0x0000000000000000000000000000000000000000000000000000000000000000"),
    .DATA_WIDTH_W("16"),
    .DATA_WIDTH_R("16")
) mem_im (
    .DI     (16'h0000),
    .ADW    (11'h000),
    .ADR    ({{11-ADDR_W{1'b0}}, raddr}),
    .CKW    (clk),
    .CKR    (clk),
    .CEW    (1'h1),
    .CER    (1'h1),
    .RE     (1'h1),
    .WE     (1'h0),
    .MASK_N (16'h0000),
    .DO     (rdata_im)
);

`endif

endmodule
